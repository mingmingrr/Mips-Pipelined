// vim: set ft=verilog:

`ifndef DELAY_GEN_I
`define DELAY_GEN_I

`include "../Util/Control.v"
`include "../Util/Array.v"

module gen #
	( parameter DELAY = 0
	, parameter RESET = 0
	)
	( `Util_Control_T(input) ctrl
	, input  in
	, output out
	);

generate
	if(DELAY <= 0)
		assign out = in;
	else begin
		reg q[DELAY-1:0];
		integer i;
		always @(posedge `Util_Control_clock(ctrl))
			if(!`Util_Control_reset(ctrl)) begin
				q[0] = in;
				for(i = 1; i < DELAY; i = i + 1)
					q[i] = q[i-1];
			end else
				`Util_Array_setAll(q, DELAY, i, RESET)
		assign out = q[DELAY-1];
	end
endgenerate

endmodule

`endif
