`ifndef MIPS_ALU_ALU_I
`define MIPS_ALU_ALU_I

`include "Util/Math.v"
`include "Mips/Alu/Func.v"
`include "Mips/Alu/Status.v"

`define Mips_Alu_alu_Data_T(T) T [DATA_W-1:0]

module Mips_Alu_alu #
	( parameter DATA_W  = 32
	)
	( `Mips_Alu_alu_Data_T (input)  data1
	, `Mips_Alu_alu_Data_T (input)  data2
	, `Mips_Alu_Func_T     (input)  func
	, `Mips_Alu_alu_Data_T (input)  reg_lo
	, `Mips_Alu_alu_Data_T (input)  reg_hi
	, `Mips_Alu_alu_Data_T (output) res_lo
	, `Mips_Alu_alu_Data_T (output) res_hi
	, `Mips_Alu_Status_T   (output) status
	);

`Util_Math_log2_expr

`Mips_Alu_alu_Data_T (wire signed) data1$  , data2$  ;
`Mips_Alu_alu_Data_T (wire signed) mul_lo$ , mul_hi$ ;
`Mips_Alu_alu_Data_T (wire)        mul_lo  , mul_hi  ;
wire [Util_Math_log2(DATA_W)-1:0] shamt;

assign data1$ = data1;
assign data2$ = data2;
assign {mul_hi, mul_lo} = data1 * data2;
assign {mul_hi$, mul_lo$} = data1$ * data2$;
assign shamt = data2[Util_Math_log2(DATA_W)-1:0];

`Mips_Alu_alu_Data_T(reg) res_lo$;
always @(*)
	case(func)
		`Mips_Alu_Func_Add  : res_lo$ =          data1   +   data2  ;
		`Mips_Alu_Func_Sub  : res_lo$ =          data1   -   data2  ;
		`Mips_Alu_Func_Sll  : res_lo$ =          data1   <<  shamt  ;
		`Mips_Alu_Func_Sra  : res_lo$ =          data1$  >>> shamt  ;
		`Mips_Alu_Func_Srl  : res_lo$ =          data1   >>  shamt  ;
		`Mips_Alu_Func_And  : res_lo$ =          data1   &   data2  ;
		`Mips_Alu_Func_Or   : res_lo$ =          data1   |   data2  ;
		`Mips_Alu_Func_Nor  : res_lo$ = ~(       data1   |   data2  );
		`Mips_Alu_Func_Xor  : res_lo$ =          data1   ^   data2  ;
		`Mips_Alu_Func_Slts : res_lo$ = DATA_W'( data1$  <   data2$ );
		`Mips_Alu_Func_Sltu : res_lo$ = DATA_W'( data1   <   data2  );
		`Mips_Alu_Func_Muls : res_lo$ =          mul_lo$ ;
		`Mips_Alu_Func_Mulu : res_lo$ =          mul_lo  ;
		`Mips_Alu_Func_Divs : res_lo$ =          data1$  /  data2$  ;
		`Mips_Alu_Func_Divu : res_lo$ =          data1   /  data2   ;
		`Mips_Alu_Func_Mtlo : res_lo$ =          data1   ;
		`Mips_Alu_Func_Mthi : res_lo$ =          data1   ;
		`Mips_Alu_Func_Mflo : res_lo$ =          reg_lo  ;
		`Mips_Alu_Func_Mfhi : res_lo$ =          reg_hi  ;
		default             : res_lo$ =          data1   ;
	endcase
assign res_lo = res_lo$;

`Mips_Alu_alu_Data_T(reg) res_hi$;
always @(*)
	case(func)
		`Mips_Alu_Func_Muls : res_hi$ = mul_hi$;
		`Mips_Alu_Func_Mulu : res_hi$ = mul_hi;
		`Mips_Alu_Func_Divs : res_hi$ = data1$ % data2$;
		`Mips_Alu_Func_Divu : res_hi$ = data1 % data2;
		`Mips_Alu_Func_Mthi : res_hi$ = data1;
		default             : res_hi$ = DATA_W'(0);
	endcase
assign res_hi = res_hi$;

assign zero = ~(|res_lo$);
assign less = data1 < data2;
assign equal = data1 == data2;
assign status = `Mips_Alu_Status_Init_Defaults;


assign \data:image/gif;base64,R0lGODlh9AEZAff/APv7mP38ufz8qZanSK+5bbjJUNKaRSs5CYmYSFdrJGV2Kuvb0ImZM////0VWFv36eZllJe3q2drpbZanNq+3jNra2urtiMfNRLvFlrqHNTVFEHiKJYaVKaq5RXiHSLrHbuvtl9eqqGtrUPHZaJBZItjbVVBlF+rsyursqMaPO+fqeLC2stnbZ6muNXWKNN3oj8zaZvjo3cnXV+rRV+zuubHGxrCRi5ypcY+ZYubsZd7nt/fvivvv59nddzNDCOnq5+33d9mmStncubiLTaq3V+74h9tld6x2MtvbycvLy9fcqd7nVs7USNSplJF0b8rNVVooHdvciN7nzf3tddqoVNSwbujtWZJsSMPLiLV7Mu73acXLqJWcNUtbIv//hO74l6xxccnNl6pzKfPNva+LcdbbSpSMiNncl+e2V///5/vqaf//94SMJ6VrKcbNZvfvlv//7///3qKtVmVyGHRME83Wmf/378zZdu/4qHlQKsfb2sbKOdvKVee2q6WtRciVlP//1uraj87XqZu2tsLJeap5Sdy5VLe8Ve/3y7a7SLt6gnuUOINUTP//zvf6aPf39+/32v//xsiXav//jMu4RLzGPMupQu/3uff3jMrKt87WuNvNyoWLNti5SM3XiLdXZoVUG2x/NUJKEtzGuqxIVzlSEXuUKO/36WyCJ/f33vf31ohsHPf359vISZyllFNZFae/wdnLZ0VUB5aZJ/f3zvf3xtGcpuSzmPf278q6Vf/35/juqbqoP5A7Sfjuufnry8yhV+i+Zc3WzEJJBgZAJ//3xt3Jd/b/jKBrM20/RPf3hPf/hJqGJt7n5Oje4tzIh3SAG/f/7/f/5/f/936Mhf/2jPf/zvf/1vrv9//3zouDGpqDN/f/3tu9wPb/xv/39//03raioLiiWjY/MdzJl//2hESWU93e5//21lVaBzdrSNfO1otfXydAEt3Fqe/39z9lOl1HEq99KVlCBcDP0Pf///f3///3/ylCCHwrOBVjOaeOH592H3V5d+/v8P///yH/C05FVFNDQVBFMi4wAwEAAAAh/wtYTVAgRGF0YVhNUDw/eHBhY2tldCBiZWdpbj0i77u/IiBpZD0iVzVNME1wQ2VoaUh6cmVTek5UY3prYzlkIj8+IDx4OnhtcG1ldGEgeG1sbnM6eD0iYWRvYmU6bnM6bWV0YS8iIHg6eG1wdGs9IkFkb2JlIFhNUCBDb3JlIDUuMy1jMDExIDY2LjE0NTY2MSwgMjAxMi8wMi8wNi0xNDo1NjoyNyAgICAgICAgIj4gPHJkZjpSREYgeG1sbnM6cmRmPSJodHRwOi8vd3d3LnczLm9yZy8xOTk5LzAyLzIyLXJkZi1zeW50YXgtbnMjIj4gPHJkZjpEZXNjcmlwdGlvbiByZGY6YWJvdXQ9IiIgeG1sbnM6eG1wPSJodHRwOi8vbnMuYWRvYmUuY29tL3hhcC8xLjAvIiB4bWxuczp4bXBNTT0iaHR0cDovL25zLmFkb2JlLmNvbS94YXAvMS4wL21tLyIgeG1sbnM6c3RSZWY9Imh0dHA6Ly9ucy5hZG9iZS5jb20veGFwLzEuMC9zVHlwZS9SZXNvdXJjZVJlZiMiIHhtcDpDcmVhdG9yVG9vbD0iQWRvYmUgUGhvdG9zaG9wIENTNiAoV2luZG93cykiIHhtcE1NOkluc3RhbmNlSUQ9InhtcC5paWQ6RUYyRjQ5QUIwODYyMTFFMzlGRTZDQ0MxNjhEMTkwRDMiIHhtcE1NOkRvY3VtZW50SUQ9InhtcC5kaWQ6RUYyRjQ5QUMwODYyMTFFMzlGRTZDQ0MxNjhEMTkwRDMiPiA8eG1wTU06RGVyaXZlZEZyb20gc3RSZWY6aW5zdGFuY2VJRD0ieG1wLmlpZDpFRjJGNDlBOTA4NjIxMUUzOUZFNkNDQzE2OEQxOTBEMyIgc3RSZWY6ZG9jdW1lbnRJRD0ieG1wLmRpZDpFRjJGNDlBQTA4NjIxMUUzOUZFNkNDQzE2OEQxOTBEMyIvPiA8L3JkZjpEZXNjcmlwdGlvbj4gPC9yZGY6UkRGPiA8L3g6eG1wbWV0YT4gPD94cGFja2V0IGVuZD0iciI/PgH//v38+/r5+Pf29fTz8vHw7+7t7Ovq6ejn5uXk4+Lh4N/e3dzb2tnY19bV1NPS0dDPzs3My8rJyMfGxcTDwsHAv769vLu6ubi3trW0s7KxsK+urayrqqmop6alpKOioaCfnp2cm5qZmJeWlZSTkpGQj46NjIuKiYiHhoWEg4KBgH9+fXx7enl4d3Z1dHNycXBvbm1sa2ppaGdmZWRjYmFgX15dXFtaWVhXVlVUU1JRUE9OTUxLSklIR0ZFRENCQUA/Pj08Ozo5ODc2NTQzMjEwLy4tLCsqKSgnJiUkIyIhIB8eHRwbGhkYFxYVFBMSERAPDg0MCwoJCAcGBQQDAgEAACH5BAUKAP8ALAAAAAD0ARkBQAj/AF/AkCABD7c0gBoFCHDJm7U40tJEnLimQYOK3yIBELBRwEJAdiyKtGhvTZxG1hpFirRQAKBvItFxBEBTQJx6Iks2kAaiSJEvXwR4rBUH4aWFSPEIwOMt2kWLcV68IHhHQg8JdxBVnPZ0TZoANCdVA3K16sA7d15wu/fU4jc4AY4tk7vsCyC2bC1uwYEAgYdFHvwiYPAB0kiR9+LgKcLCzRM3Bdx8kHyG21M7gI5ynAIkRwcXLkKFDiVaNCciRAocKkCgQOrUBT5gUWWxokVEFiSoyKFCRYC3LD169AYHJsw1UvqFErG8uQgEPY5xBvLgwbJlyggShAGjgynSChSo/1OQQIGIG6wOPzpcb40SCSyWxC8hwQKAL/cDxGnAdo0OcR0MEGAHfnRAxAtBCYWHHAkk0IWDXXRhwoOhaGJbA+tZtB5XOCFBwAQDgCgiEUqIhFM9cJzBwkASaEEdAC/x9xRXp5yggw5KCLJFHTtiIEVFukSCBxArQsaFAhGO04UoXSjpQBc3ONUAVz9QwMBgDFyJABdynGBRBCiAAEIPMlxwQQuzZLkIA2ty4sErpYwjipxyipIAAUWAgAgi1kByDSsnNXIJIQMMgEChISJKwCm1NaALWDTV5NKFI6FoDUuYLhRJGhfKFOkxMMLUaAPcTKWbBD4d80UA3gQAlFJ4BP8AqzdpNGDPRYoVIVVVaXlyCaVQCeDFsA9oAcOKK3IHwx3WHGYRHAIsQ511ADRSUYYNYIAAJ4uA5u0ii2CBi0gX3pPKF0DAUEABT1Sy7hMFwECDSHA0IhwmOWghQQeohKKAv+EFjIqAHXRQgIEdHJKwwQXMKyNbvuyWw8Q5CGDHGta0qik6tnG1BgYikOdgg3MkIMcXmIwwsRU5OAJEutxJsIQEhzAAWngNNpgHDhE0gJOG7EXzAgslLHFsGfTdl99+JAmBxdNQh1HHHfZxJAAIA0gYYSkOdP1kP1KMhO16JzYghBxcTMAAFwxMwKUSwEajAwgWqMDCxECsuh9eIgn/Q8QAcgAOuBxy1CFlNNZ8UYR2MEyASgImdC2KKBpMDg8Ftt2Ki5VscsAGB5wwIEfPa/yCwgsW9MCEmS0w8DkbpmzAxgbQOKDBAbfn7oMDcljwQg/KvnAJIN4I+QECEywyGAKLGDoAAek1AJNM1XhxzCSRRgKHs1PGsdBRSAXQyPYiPbpRpNY6G40SdwzE4lRf4IFHWgjGP+v2tqVxyX2L/85CVhx6SmLwcAxMXEcLMlCWArMyqmddQloPoE4RvAGTvDyCAB4ATWm85QHDIQYx3ngZC9almhIewg3zYosdhCQUfOmrEv3CGXlmiIoJFMxgHUjEwoiQw0QEghY0UEIg/84QiB70ZgoW2MEUyrGDciijGspgIiZ2YIFAgCAQKDgDAbSxgTmUrEH/qsMlGLOEMi6BZTmAV7wSWIDkdcsFMkyAB5AgI+75bA2qkJ8AdoGHXQAABEDJT0jYggssTOCQiDxkB1RAk6C8AAGvmFAXvNa1LnjAMCLhikU0aasGaGIAbVtb27hABB2QyyLSiIIMmMBKVpagYtfopEhOQQDnFQoHhfrAj1ToDcW9jCAdWAQqHgchyYVCGCJZzyMwoCbPgU50iLBIDFBggdQ9YQ8XqEQLXje72dXOB7gLpwY0wDupwMANMJBBD4bXKjwQYE3giie4cPCB6FmkGABQhheso/8MUEVCF7b5WQOiAQihGDQAHgFEQE0SCaGgLy8jWV86YfABGchAAjAAwjGKsK4PoEUqQGnKHdcAh2wgVABfOAYQfNestkjPGkVwmSO0gEAZuMGi3EFLNJ0FBzxgAgjKACoQArA9UZ3iBqEJDSoU0C9UeEAQnLzQGmphASIdrBI5NBgRCJFChhoUABOTQAGWGkfxKGAOCOjAE1TghXJ4oRqTKIdY4vpWusrVrXg9Bl7b6gV93vWtfM2rW5WxjMEWtq/lqMYDRsCHJ7AgFzpclwza6II3atBfHtDEYW61yTuigGglCC3SWFAEPAjyKbggRNqQ1zZFqgBlbwCABDihtUn/VjJCOGBUJkUiKhl9cm0cYEBwGVDKD+5Elay8QCtZ8AVa2KYi9cCAB9wELuYVSglcwYs1QAAECfyyA2zyiwc8IB4H3aAZT7nVI7BwKE6Ygg0M4AQH5LDTaVoABKosQCWwyoH3dpN26bjdAQ4AznE6YABSmSxk1mmNo4BAHNziYGUDgwEp1WMaDwSCyyL4AAAEIBW26U8D7HCJlOLnfAEAxGG4wZKTTkp9Z5CMggsggw94FwgBGgBqPuDRO+BBGhiqyBrQoZKT0gQPnPIZubxRhJcBQQtpXBdkIENRFJBvJGu4xJOf7CKiyvIUOCANwP4VCqcKwVnXwoMKtDDCGxZM/4cf8NJFUiGrFlJMBhsIDzRaoIJlPMCvfS3sMQBdDr321dDVAIABCVvoKGJi0IbuZ6MFzehBH5bRgR6sE7FTWE6XI7EA2MEhNgAaTngrNB7AALByouQT9CC0MiiDDErAgrx9YRcBCIlFqpS2UCKSCBb4CSDvAA1Z2JZrT5JQlCyCE2zdaitrEAQosyTcLBX3MKyIwhOesDomcJsFILgEHCCKBA+UZzwKcMFfFmURtjyil4pbxuLUBq5Tg+cD7xAghjAgX9j5mwN+kLPp7ksmM+13FmxIOKlp94rbgbMdBN4dDhIcmwL4OBJHeYEcNOgCVCS1sqp2SzTw4LKXydTDqv94bm1YwY1rxCEVgIB5KoriUha3BKExGpU0PDFlElKZpt6BZ6FQ4wlMWiQN2UCJQlrsXKDVJoRAUAOUVYCqVV3j6txIxTU21JapKkPqNM3BJUKSISl4AGDlCVgoPGBKcq0BSHiQQA7a7ObImvIeQw7ALhQ0sRLwQQUPKMefsWNpww7WC1NQwRL3OlhQRQoAk3i0YNsa6U5j+vKXvvQ+2xp4zu8Vro/Phc0AwwkKkK9sznJ1rGPNhDJk1LRvqIWuG3ACArBWbbj/wBd6Emw3KEAUDhBFnEqB7ARgzmfKZDVJpoEBtlXbFFkiwI8E6ihtK9dMF3gCDCzgizSIKho3ODb/PB6kAE5sYQ0CTQUKtEMQGbCp3qd2AScEceX12CMMgwHXBhYBOxzIGUyoQyaVsAf7lQgG2ANKIARKoAQIcDsQN2DgJAqcIAEv4BrrAgMvICsB8AJh1lRMRWaLcH7QJQ27AGUm6CKrogrkw1nugRYEoQLBVlqWcSFBEgAtph9C1hZpUAeQ8QGrsS6HcFE4tgHD5HEuMAEIQABtdxFpsBJOiCngkDmXEQBNJnU5sATrgkM85BqekAqHwRbegAmc4SI5gAdbYRFCoBw4A0bl4QFhk0wikQogsARzVwAtMCAFkjBnsAZ4lw1LcTWxMALlMAUPMAXKsERLpAx/9mnlwAIj/xAMlCCI5eBp2FEOmIBYk8honKaIUURYnbiInLhpnViJgveJnehEqHiKyrCKy4AJkmKDKIADnEAAqVA2q9YAEaA6ZdBKsqYCgBR7vbUAciBKzscAA0AIu1cEwZYLcwB8k1M5wOcACRByMjI2U2IRJ3ADzoNLXDAAOCAHZ1ZBFhEN1rc6F4BN27cL3mcRSJAAw6ABpeADkxMhA2AYEBUBQ4NRRkMEpmAKHvePoBEYP7IGMEE2QhAiwsUG/GcKCNB2J3A6KgA8++UuaCI7G0CE0GACAnYAD4g7HtADFYhDHxAIDBEAnoAAZRYw4UEa5sdb1mABU5cv3hUUTSc9FsEKnv/wAfHyATFTEFIShwgVlDZRERB1D9xwBpOlkwdzMG4gAVaQCNCgdqLhAggQBh0TBweFFP9kG+tREXABACo1UzlwMG6GMFjghcchI6rwU05WMbWiIVKAARRAAB9AADdwA3ZJABTwI6zGFr9gNzlQAnbYATZUIALiCV5JC3gQiIg4iIV4iIX4mIY4ApQADCNAiImYiqD4Z5zJiaCIioJHiKXYmaQpeJ+GiDMgiISoiI2JmY7Jmp/WeYkGAD1AACdwIQJ1IamgSrvIShbli7eWDRdyNtRWbYfiCXhANxbwBgRgAs9IOeNUCnaCAR9kjSdCS/HVX/0VfXLWFrhQB09gJtj/lH0woAIowDSPcAPjNE64A49dgAHUtwYCwR0JJAN+ABrDVGb66QI3AAlRNSUkBQfRAAfSEA0DGg1rsB4RcEUWEAUlUAkXQAn71QIL13EbYALgNGADBnE+IAJpoTAFcwg98IfGwAlzQB4lY1YK4AFbwFu1IHcUkwPepRTOdS0WAQkUcAirwTAJZIYuRWcGJRRx8J8NEBUUBRlX1QFNaQUFsAHl8aQBEyXNRoWvKACRoFAN9A0FxREqBQTtUjAFYpiEEE0QZRGqUARqsGVTAAD7IWQgAzkj8yANggA7BSyuVjQyUAkT4AcD4Ad+6gdyQACG4R4sEAhTcKiImqiSOYhq/2AIMxAIh3iIjtmaTlSIg3ippxkIwRAMVJALiBiZhzoDfKCag/iIhkAFaGAJnSCIIzACajCIM0AFVWAAkiAOwTACkrmoi8eIPUADvYUtF8IKAlEC3NZK9ZEn1tAf0TZtwQV9onMGyQkCqCMHrzAO4zBOPjBOlJMH1NluGAKHHHJU8ZWdocMBhXGNP4MLD0k3RAMDtOaL11ARmSAC2doOuVM5IvCGGcIDhEBCNBZM+WkOYiZmN6BbFcFZJ5CFhNkCiIRduHg6DfpYBFgJEho7F4kKGZmtk0M5w/cKH/ACOIIjL3AGgXQIUUkeIgClzEGNrIACE3M3dMgCU7B3tUA+ef8hBTwkBwWzhR/wK11BKlbTEeNjIlDxAu0zWQWQCEwpd03aICYAp234f1HAIj5RE96gcrWBEAqBULIFLyBqmIfQnd6aChZAh/mSA5iwNz5DAQ1SW1qTADhgdFhGA6+2BHk6C0/gqq6qAmrAt3yrBlMAuIoHuInKGYgKBFMwA61wqJC5RBYQC5Y5iMGABmgQDFVwqmhQBVQwBE1QBVVgDA+gBqaKqlWABqRruqdaBUOQAkMgCbJKBamLqlQADJxrC38gCZJQCJbJuIdKmQYwA5hZiFMQC4EwBr8QA+DAA6nwC+AwSNLDQnwEAiowAirwAmLCNAkqBGGAAVjwAXKJAd7/qwSXgDovEAWHoJcfwBcKqTwIoEt8+HbfCjSaBAk3EF8LaQocwAGEkB44MQ0VkQrkgH0Qio6+mHKn4ARdsJ73Og7UICWchQRy0AIEkwiOo5Jp5y+hQI0Hi42EgKQ4VDA6gBOqQE341QMFsAcSul8TMDsbEAoZq6EwrAF5QAgvQJh8mjCA9AXiMAdPqzUT0iCh0KIWIYfxER9lxALLCQA1qV5KoLM2tKcFUgA7NRKqQBOOBwCbchhesX7cQWNZuKSVkJFw2sMJIAJbwBUn8AGwwR0w+AVXixMXghmNsLVC8QUqkE5JWzDPc3cfpAoqYEYyOkGIwbYO8goR0gWGnAA3/wBkcHgRZ1ACZSBregpKhzQL2pACuTC9fZt4M/AEmyy4gZuoWhC4huC5gWAMVdAEt4C7VEAFBmAArXsLfRACs9wHtou7iiAJrbvLuNsEqizLshwCq4y7VYC7rSsJt0DLytwHzBwCCxADYyAJmosGKZACBqC5sHuZiBoLlgC7VWC5z8ADMvINBNkA0LIb80GsLOCL5ykSrGB78hXP+WubtUA3U8EJpaDA7TlOCaBZJKFkncUhPyAHsxBc+fs5DIAFyWcbrBAGF1AA2USAF1CeZ1ALa7AC8TAOHClOBxAKC3BKuMBvWYJ7FwoPUDtDKyoI7HERJ9DBWZi0rqED/3sJb//wBXVzTZSQCxM6C9CAkRgKwxoqwx8QBQu7p4cAAjXtB5ATOZPE1F0QCir9JSpQNKEVWkj8BnggbiOBC2HQpxPAsIXiB4SQCiJmEbQAAIV2PR6mC243DXHAxSVgUeySCBiYAzKwCD0cIYZsAmbMFQtQSx1wh0oqAy9gj1iGC0tngzYoAJhQN118MIewh2LTAKkgEEQjHypACyLxDjfQtpLkAIl8A+RDKdIQCCXABKetpxNgCmzDBeIQC7caDDOwqVQQBIVwC1UQC2oQCKdKBa2aeEiUeLEwBrrgDGOwADwQDowABXkwBKBAB1DA3M1NBmSwArjwCLiADXbAA3aAC3b/oAvf3d24wAq4wAMLEALdgN590ARgMA5QcAVXEA/MjQPicAXhgA3T8A7+AAbs0ATrDQyt3MpBMAKBMANB4Mq3Ggit6rmq3ATukB6PAL+PUAtPdrZLUAYSAAK7sAtrsWv1K1+LADr5Wxi0YL2/4wLQaa/i5AMKEDZlehialI1cYND9tSZW+bMNwNXZFNEQWp7CEwEeEE4cijui0K2NggQD4G/+FTnjcFtPqwA7EzbkbKO0p5T6VUINAyQntQsWAAPnOLEtQKG0Aw3NCNQDpgEJQAhRQJZGHWxAMACfTUkR4gFnho2vFtdIQ2vLmdUr2AA/8AGFIiKIQgiMfCG4YYhA/9CKXkaU5gwIIIBR6TRZk1WeWrAEE2ACTO01ExJywijoNtQBDIR6RZopSKEgyfkFu3IHdWBPqPUCsQDJcd0DviASP4ADPezUP0wBmzXEd7CLq5QLXDDjWcI2ICLT2RAFbsACoiu6sVAIuiwJAA7gB24I1Mvs5DAGfXDcCzAG3D4G64DcukDePBDuuFDu3i3u413e6c4D667u3M0K3R3vPGDe297t2g4O5CAO0l7bs+vK+7APBoAM8bCxoUBHbgGHQlYMO+AIU6AFVjB1WN19IhEB9ZtwCilf+ssKqoA68BEK6ynkuOMDocDHnRXQPiMFoNSs48oFnsBJIoEL5KBfEf+6X3sQC9VLAxTQBeF05h4ZPXnBA5ogCHWQI57wNw2XreTEJHJasKeUIRGgkzi0lAUg0w3ACi3GEVOdXNlECVrCFzpv5hrQBYQQCGJFloeQREUASV3T5MCHbB7w0RaxACyA2q0XayywAzXtC1dmNmjjNkh4SANwBnDgMSJxAjIzMS5iMfomDY4OPOdkU5NeVTlABCXzJF1TChFCAVxBnLjXWoRgGP0rEoAglEHJtRsVVN0FkmkAxzKiCyDwBBa1iyzgMA1gdoc8SREyIQqgwbKECLHQSmaiNtA3XMEON7QAArGQC8vuqoZgCQYwu0FgAMBQzRmQBUdAAoXQBNJMAQv/oAu6wAOsAP7iX97h7+7mz+7o7+7bndyjYAfbXd7fD//sDu+s8P26AA7RDAzRPgTbABAGgFEBZmiEGkqrRA07oGFcghoNJD6S2IDimgb3aFnQYkXLxxxAAAQoBueeRCk4GLBh48IUm0WcwkRL9QJEIDdzfGjQ0PCAj3YafIQS0sBevWkN6lVcivERK0iQIkiVegoSLooS12DERe5CpUqU9lTaE0tFlCiherY70LZnl0wZ5TY4McDUBhcbNqCao4Gtj4YaRJXq0oVCtIoYK0IidKhDgQ6JHh/SkVRXpAABBAjYkWPGkjJMxs66u0GBg7ap27brQihQEQkSYMiAsfkL/4JXshyMEzVYlAMHHqRIhHNGBhPkyMuwsADiiy/ERteEGcDA+gQG2OXoSFzxRI8yJUosyfFFV+I1cSK9YHHHvac78D0FUpajgIIEhYETdoDjVANBqsPuOgQI+U8rrWoBAAABGBQgswC+OKYIZSi0AAgU0qioAYy+QYEPGZ4oQUQajGpAk1CA+20c4ApTAAPFlmqKBjf4uICJCwrAzhQGOLCOAQTq0KWWm3KZ4aAZDDHAEoEMCKLJJ4FxUiAqhrhiDB6yZIWHLbfEhUsevhQTzDG/9DJLXWLIZAEyw3TTzDd50IXLGMhAhoopqQjCkGDUGIGXeXbqiacuXKnoIhMVg/+khyVGyCEHLUIaKRvFGhBCJZhcaIkTBJRYQxcdXnjBjQR6Wi21nqCpAw6JljopqaUqyoSTRVzgxCVOGODCUw5NbKCrAsAStpInJOhBjmFMRRUK/+RKao1NEGBDL1T2MgGo1NjiSZQutpCx16wYc2xcIgogQglpGtClkcw2A6AIFSxQQQUWWHBjApZQeUW11HxIBgsQAPgCE3glyAwPBExwoJTeBGNRFGqakYgVT5jgA0ccZejBguZ2YXUiCrj40ToEGCDghO4kiuAOJo4rQwYQzsNoGjgAWU8GN2QoQGedYVBBGStk2CC/LvZzQBYcIlgDA5F/5ACBAg+cC45dgAD/YpkHJmFQsyKKAMJrsPHQsFd7JKqFhRLKCA1mxTIRoTfeNGC4aAXCUAyjDlGI5Ykbc5yAA044WARw6whR5RILojByhBksQWOEEZhs0oAmpbR8SimfNEASSa4gY5Qss0wFzC5JN7101E9nhZUY7FhAEkaGkOTyJ2t3sk/I95nnJ594GoaapHp1akNVejhOvBzIwyQAQBS7R4kBuOCAAzZeWoQLHdaIhgYUXvjAhLUOYEtbDbQh5Bq851K/gS044QQv+DngQohK7VnjnkdO6B6EHliIRYZYRMENClANMdrigy4UhSm/wgBL8lKtUOyLLarRVhc0saFKNQASBCBCBzrg/wcPSkYJiFFPuxoEhBxYYQkqXIK9rMMGExwACvxyCAVQsKAFHeML3ohDLW6AHxOUgmGlkJsokhYHXdBIBn3D2Maak6GTaPAGDODRIkZGiFRsyDt3eALGnhAFVVgkI2nIRiTO4IYCoLEAO9uZBZahhSVwYA4mUFgXSnG0UCABFwSgYo+c9oEsTkQip4hCveaVNQepAAiKvJAiQdC8XiXlG7VQQQ7QJgMZvGBsK+jCMEQhmFckQDeiCIUmMngRFHSxb5VowSEogAUMwBILWHDHAsghjhGUgHG7NIQ4UmCAX6ZAHBg4BS6w8oh3PEKZ73jHKU5RgSRQwBXUwAEZyKCIEP/YIptNaEII/kAGMJDBBiFgU+h4EAM0xWATNnACKWRnOWBcjnaVa5IlggA5NcxgFvPoCWDGx5N+QAJBWmzAN1iBAhAklGM5UAEmBACIxGjCD9Fr2vQGgDI7hCoKBHgFYPgVGDYUAAXfcFZFgqeU9k1LL3hhA/YqlRVWkOMJBfiKsPjQAy6I4qMNMUPwotiACNxAL9DYywbmgJoJZusnIhhOrwa6wQ92YAJR7cAZWLEGmz3IXZGyQldXqIIXyAE7fRmU+AJzgxMIDIdfCAAcUsFHVChAHQorxTgYxokeYMICPbjABfbwlb6WYGM2scAb3vCFvYpscIPLFQM8ER1f0SX/Fn17wh5YQIs1TGMNj6gFHgTQA8iEdo0FgAEIMNERLswBHnW8owNEsIWgMiBw02vsBwSawV/EgglPUBt5gPAFEMCgXrFRgQTAag1YNSB41vjCMlDIgiW8IA4YocArXoGARFDCErngxSqG4QEFVqRsrACBeJDjN+pRjyVsYAYlYjGDMsygBDOYQStScN/7GmAI+gVmOITxjmbogR4CJvCADayHFVTAHxVYwCi6qU0INyHCE86mItixgiToQcMHPvAKzDA7yoU4xL80AJ8gN4N9rGInSm1HO3ygjqbeox6xmksqjHEBSgB2D0yIggDQcTdBgHACQ8YOF+SAsjXQ4AU9/yCCLDxKQw1wQqQfE6MgJ4IBTrCBqHjR1EU3BNNn8K2vgH0CqZ58qm4tUCKZQICmiErUORTGBKHMwxxCgQMz3IACPxioUzc4gAn4IdAt+KAnLhGAS2xG0QDgagrJkwNl6IgDGxCBAkyQHxF4AAcIEEcPjvFpABxjeW6lQHXaHNf8vKILCIgCJnbAgr5WArAXKEEULPACCwTiDTt4gwXcQNuXmCJwXGCBYd+wC2O/oQd8+Kus91ACFfDa1TsorBsELVUPFiART7CAF4CghRbMIQEm0E/RunADEPihj4ELHAOwwAotJlnMfENODjChglyskTbGik0t0gerNABgElibgv8W3hCHjLjiClzQbsMp8fBccIECqdjKVhrAihfAIG1laAUTWjALlmgjEcHgQyvqO4OS33cIKVh5y1OQBWTkgxFOaMIWFrCAGEQgBuiMAA8iUAE9KlOZuHDGJvzBc3/wwB1OGMMCxhACCW/TFjbAZgicAc0fROMRzaiBM2IAiRiAY+cLCIETrsCIKxRCEpT7JTDoa4UZ8EIbChjGk8OnAQsi6CQ//RU5crGPVhykFZVgwRe40St/EGIAUhW0oCdAgNv+AgRRkMMqQlFpEYRi3OkwQTo40YEowHt4fX4ElrVc1FCwYQAR2FAUuzJmZ1/gCVxY8al64gE+S4Ska1AFAVT/SlRUQONa/ErqMBCwA15bAPm78MV0ESEHLnBhAtIP9ABg4CBFuwsII1hC97m/hAf0QKoK8M0nt+UDBKhgQsvAxDKKEIA0/HkAA1hErVygAPzIYUGv7muz+8oCXAuEXEO+NwiEQ5ie6mGD9OKCjSFA5VO+HngCWaOEYJGBaEs+ebEASZu+CSC0x5AAZeiIFmAAF3ABVHCBUEDBUEAAGPAD0qAiDjAFH3EDC9iFMxgCBNgGCniBXAAssqC14uKFFvCDQ9i2J4ABGEABKiubegi4SfACLygHLwAAhLsHG0iAVUCGVeACXmi4Lnw4SsgFMeSCZ9iFEeCDEpCBEuCDRGgB/z5AQz44OUPghW3IgCywwwwgASfYhJuLgAXwQ0D0Op37gZyLAULsuZ9LAn/ACmwYOmEQBkLchFFYgSawARswAydwAjBgOi5ZgHBYgXMKRZ6rgEwoJmWSghroOZ9bRZ1DxCyJAbPLhRFAA2aQBWVJqhrqEImwAwyoAmNQAV2CHF2irxZIhFhAgSzCiAggACIbssbDgnRpAFXAgyhAAJ4wK1wUBQZIhDtAhEP5RpDJspXCC064AW8Ex5gKFh+8gBbYF2U5oFf4gHgprAfsAZCjlr2Ahi54R355BXHYgSmgNuQTyB1QAenxEQaYheyYADf4guxbtFfrvkZpFCDAhCeYgP8NGKW6GiJR4AILmJCu6RoBSIMTuIEBQAD6Q4D6qz8XIAQ8iBAJ6CL/u4AeeAEVEEDl2wFMiIUP8gNC44VE8INEOARbE8gH3IEIlDWlZIIcGEiOsckCmAUfQcgh6wAYAAIrcIQOELf8IDd46AIT4IQ7EDQemR4Z5II7UIEpmAJKYAZe2Ie3jEu43Adt0AYXjL6qfIwCiIJaiANASANdSANuiAQAgMIonEKEY4UrfAVkaIPGhADIXAUI4Ich6EJLeLhOoIRWeEsjicP5CoZgSIEM2Ac8LIQsuENkAAVJWAAGu7kFcIY/jE1AjM1CvLkYWIBMaAZ/eARsMCZcwAZnSIL/H9A5nmPFVUSn4nRFV+Q5Z6iBZsCKZJKCTKiALAkHJ8A5Q8w5PzSDK6AcPuGFV9ApDRiGOeCCWIiFXRpG+solxrGvFOAHhsuFY4Q3iVgAOciO7KA+P6iDaViKVBAAC+ACTzIrU3mFUMgDLkgEN0AZK6uyBvAHCsgVB3KfcmS9ioiimAKLYBEWaEiWuxOMbZAXo9yBEfADbZiW34MGW9yptkgAQgCCgAQBpwRIg5yWl5gekSkAh8Q+BgEAIICu8QhSFQCAHsCXURIFu/oNI3oDsPkaILgEaZACk1wElaxSKkWAMwAEQAiAZUge8eCbJziLm8w1EFC+WOCC6tmALDMF/xfgACLgmBmFQAn8ij2gBKYcSAEMBBWIhTtwgzuAgf5RgR4oruSxggIQvgRYLbAES06AAanCzz5iwIFEPmPgB1DIg0vNVEzNg1VYhdHkBV6whC7shBlAz4MYgUBgAT4guTjkAxbQNWTDAQXIgwR4hTwgAWSITAiQTMkkgVXYBsykhE7oBPvKgG0YgkLIAGVV1jvchtPMAtNEhjxYzZtDAtd8TdmUTWfwQ2dwAnbwr0XszUZsRH8Qhk0IxZ5DTnSNAdjshqZj19t0hqYbgzFw1z7ohj4IARuwBVvoBnfthj9wgj/AuVbcuRiwgStwuRTgBTRAOVClrxmgAkvIANEcgv8MsFhm5YdEAItEyIUnQAE7kAtNwAF2s47o8wNPOQldCIBAeEs0zCX5MoRVmId08IMcOwPFoAhXUa4GaAY5cKCWYIlFkIPb2go4SANaoBGwyIWNZSVbDIreOYA5cINpQz4I9IMN+L29QAWdIj6fwKu13IFAGNGCbIH1yloFZIM3BYA3AAA8WJAGKQIgXYIgVYN3SQQ2UBGOdICOfAMgkIBFAoIXwIM40AEcmAAqTdwqHQDpioMAKEznsqR64ZhbyzU4jThOeImWeAkGyIVJHdERmNNKCBYmGAFq67UMdAOQCzaYYINZqIQlkIEyqAR9zA/b7YIECIUP+KBmlB8/UIH/N3C1N5BRYIy4dKADTO0FUMiHTGXe5CUBEoDMI0jWLGA5EZMSKqACQ0AD0ByBYNgl0DQEQ7AE8mUSXrBYfuAHCNDCNnDMNjgC+D2C08TDO6zfDDBNeYBWZEiGJmi6a8XWPszWCPC6BQCDXjCCTzACBV7gBf4EMGCHT3BgBwYDRVAEbfoDdgADUtjgCP4ERfiDDkbgT7AFZ4DNTeiGcPgDM3jgT+gFM9iEH9jW2DyBTTA7i61Yis0Ax5kBNLAEZljWQkAGSQAVNwjD0a0Ej0UBeLuH6UCALNMGZtgHSojDGfATP5mBTtCcX6KCXFAAWfikV/CD0b0Da9gKXyjTXtsF/zX2hAFgiZVCUV5IKF/whV0YW3mplxJAmxHhhBUblKAYBjnYgWrgNavdATdA02nJiw2AhjlgCGxEFVEYgCiYgqNUvgvEKamULRzlhAFgAb36gjfAg7b9gi94FFN+FDXABACAAS5QGN8Qoi4YBwSwgNh4AQmAjS+4BsO10ioFkgHQgThw3AYJtWOwGpEg5eagXAs4QFpZr5cYgFgoSDwdyAjsqxzLhZsSSAHENULgAlpxiQTkgEQogRuphIyUM9xNgNx1jA5YvAkAtKnSyWoIXuRTARm45q94gkRYhXjIVDrw50slgVvF1fetX+vdr19CaP5K6IothCNo3+iNaOiFgP+Ihsz2FYP3lV/TvEPqtcNn1egsEGhy4sP/hc0A9sPbHGBYNIMYwAZ/eOl38IeYjmlc2E2bfoTddAZFSGAFHmFy5U3efIcVAAMH7gaXdumYfmke+IFNyIRuEAEz6AaTXoBuyMQ8mF/75Wg7TAFgCAbx7QQ0+GpD6ARDoALtsoT72od94Ad5EAN5cFb5lV/7zeH74gUq2IZ44NveEAUF6ABZuwAJqOQRjQV8mbSgVUBeEFHls2MVeIJcOOJK4IJ0iNptWYUeUAZMoGe9moJDWIlbaQkTJCuf0Jag6AIiiDbBRm0V8APNzdoNoB4/6IFeK1NqA2W5FQ8WgAG6hTQAsAD/P3Dl3ZgbB+AEC0DCWpaAL7AGJdg0xVXcG6CBNBBmHFqQSRAAzEA0ANgFtvVtTa4eCY1tsR1RCIyFHuxB2XOim7g1FejmwIEJxmKAQygBpdQGWTA3ByiMBFAAOXADN/iA/naDQ/iAXBhSthXeQJCB8sax846CFzgELtiGK4iHebDVf/7ngYZMfkCG/B2C6nW5/Vo5hl6503To9oXMij5xi4aAi24DMYjr+c1fjobWLNBoEmCETOBDay3pBZACAca5TTADV+ABfzhqm65pnDbyRSzyJEfymm5ybCDyl47ypPvxFUjpbP3fmxsDMLjq/M1f+fXy+G1xMX9oMn9fFjfz/xXHaIw+ghaP3yz4hFV4hRYhjN8AjlCgqSd4ghFYbKOE0zNtb+thA/iG00q2AL7pQbBAhboaFJ7QgFcI5OB9g3me59X2ZsCplSxTgEZndJ54iDs4yrFFPsb2A8Chnhtlg9guwFsr0zK1gEsSD/FYgh1okJxokd/gD04IhA8IcBhwjxe4BEHAgZPs5ZMcAAJAhDQABHcZZgaJBL8EhGLAjAbxbZFxYpNlgAKgR20e3gKcrJniGxnQtYQKhJsAAcWzDiuyDvk5BBZA9FlQkS7glnRehMjogHHpgHJxyAYRgLa15zwvAMeWvbPwHm9mACvKFU7gAkKwAHFYBTogAVCw6P+MPk0Ov2EPZ7kUMIIhMIL7PQJkyFWKDnkUj14VV/H3bXMZj/HT/PIZLwS064YFsFaZx/KT/kNnsM4xcIYscWl/WIdwEAERoIZM+IGXbvIhP3oiT/qjL3oP24TZnM2bM+lNCIFkAINxWgEygAIS+AT4zYIxRwYxaHEzx+jGJPszb99cbd82WN/1zUItZAZdewNCWIX7bi1zA0sEOI4QkQBC3rVeI0DC9pHAYSwucIMdAAFuL6wytZFYa4F0QNJPIiKG8YC8Sra2VbboQ3dNZgBN/yTzcxhSigJeQ3zENyzEpzZe0OTBly05kO3msAly5xgWkAE0FJE8toBp9wByk/P/FukCBbgDIpCDQ0ijD+iBXagDYUdJlBR2YT/2ZH/IzWAewAxmv2yESEABAhCr6uAClFT4wrJ8YwsEGHiCEMlzGIiC4S13cjcGOUAAkXl/lDyECJypAVC1+x4H/O4CFxgAIgAIIocIFBB4R4CAAAkRqmDxRMYTN0+exFIRCIQxPwwQbGTAhcGEXCDekCSJqQeMEiNYxBK3bdW2LENk0hxiJIXMDDMzFMrSRgyENiQgDCVhlCjSoRCQtWl6REyWnkeyUO0pL8vUI1pJMHK3aQGSBWMWkC1rNkJZIex6JSNwwxw8ETa6LYjhLEYEu3j1xojxQ++YTYJXdFsRIpwrG4lt/zA249iGGVcrbCQrFG7UJiSZhWgexY6EVmRH2oxmKqYNU6ZtgkJovdp1awig4sHkguBQoDcjSRJS0KWLg9/CuyQYUKIESwlvAJTcRXKksQEeO3IcQKjkc5IWYk18koiNAwfjHIgSH5zA7l3pA33gMgDBR44IBhCoL0cOgkWcFnngxKXHDroJmN0bOxxiW3weIUBEFLqBcNFFL4DA0kMPwcCCCgAAYAEOoSiggAgfgujBB0QMQAQRBRzixgtYzIfDADjcMIAcN8jxASJpAIIQjwhFEgccugQJRxxpcFOLDl+ccYYnnhBiDCGegOAclVOSFEgPbsDgRixu3NEgCChcBP8CCJ4Q4d587g0wQC49UPREB3MM91sCXYSyYAf1fVDABy8E8GcAkShkgQQssAADDHzIEIsFZ4Ag4ZhkgmDBpGSqR2UUMMSCXA8sfCEAIf15MCononJywy4B7PJMFUMg1RooRxk1q6yvwsaUVlplEdNVWclzxK9ZIJOHDQtkFhayYJlFlhAiwKOOOfqIoIgt3ei1QAR3YesMWtl2yy224XZbFlpSmBUWWRUYi8QYmrkr2CZCbEJBHlf8hExqTaG21Cok0LHKKuJUEUhub0ThxwBo4uAeFx+MlB4BvtWZB3F5JJCAAn4YWqgKb/CIhwBvUGmMHGhOkKYfhFwq8pQoYMT/nRt++DZnFyaE0kNzIr/xRQ9nJrzmzwjUKVxwwRGHQBQtO0cSlSTlEnTQDDpIpoQSouSGDFjH8qWGIAh9MXEXwxNKfTegWB8hdRCwDQ4w4lAjETcQgAEkOgJ6dyNprBENHHzjQiQiZ7xwhycffEDAIVVMKcAuvuyCxy6R4wFCFFvHwlIPgeyCAh4oeI7CGR/cN7o4931Q+R1ufHDDDW/L/XrbZxNgOCEveGNNJNY08ucuFvSgQhRR9NBDFJ+fQcDoycuB3uPN44FlLD1E//sbBIzqAQIevATwNj1lwRP4PUl1BL6tFUVrrbGthqtoU0kVFVZPxX9EIfmQ0e5XyYal/666C2SSDDECSIwDDPAAZtiEM8JlrG7YgAxmYEw3NhGDBSSwghQsi7nKoq6w5G9dmdlEYDSzCcyMYhRmIMEVkEGCVRxhYE2zgJZioSlNqcBKUSgdjYB2nzugwDmQ20XEEiCCiwlRiAoIhTiGpwLqKaSJu2DcG6pQBcSJgwBVrKIxfug8l6GkSx4gYtgupgAC+NB5m6uCHPyQxtHRCAEKgAcYwRgKIvTAAmWEnBZ3QQhx0OhtOWTQF8LkuTBNKRCpm+HWehC5L9xARBgLkQhCsTwi1AdtnrBe21rHOj3V4RppiEMkQinKH8Fhb2uYBhxKKY1acM5zL3hBHTxxBkA9sf+WknuQJ6LwJeIFAg80oAEKfomH0NWHkpUkQO0C8YIoeCJ7IvBAJJ/5TBy4RU8fwAIKIlGLSHgDEKpoBB6+QCkLWCAKEtrcLpSAhWK65Wwf6OElGreLS5xBeFF4hvBecDzsYQ8BbVsTAchhjTjE4RoEjUMjItEj3TzjGeIYwirmQAc6vGKiFM1DHkCR0TysgqMoXAUEQCrSK6xQBFeI5DYE8Usd4MAJgTGWsr6ywbKgK4FlmUw/crqCGtQAFj39KSyCKtShBnUQsDDqIFYwCDN4wCXaWAVJQ8qPFFIVX1bFF2rKh4ylcDWqIQXFKtLxryqAThxEWJ7Z5EaAM9QSjwT/OGkoohnXUISCEwR4QQ+WKaG7BeASfxIAOQhASTmc9axrxeM85+mLyb2APR6YqzpAFNcbBIJxjmMc5FBgH+QZVg4U6JBcIRlXBBDCIpdNbDzj2TmXoeAFrCVk54ApW84FQng9MEYP7kA8yYnjsdCMKzQ9cANCUIC4hMAAFurwWU3ewBWuoAAFMKCEIn0yDoCwbhy4kQY4NGAN3W3APdZgtz954xKX+OUlrAuIYkSiGAHwxXtVBToQCE5wKLiEL3xxAl/Q4BJKCENxA4yB4oaBvvWMQus8gAMFM1hGH6DAg4nrCRq0txHWAEQqAFGLvr53tfClRS1ocIboQpgAFEAm/zYX2zhfXAJ09V0SfTGpYLexjgICJagu4pBjdAhKUHeLBIjPEAYsYCHAxD1DME9AAxZDNwnCEMY61lGBCpyjAs2wspWFcdRBuGIQXnauCMLcD2pQY8xeRupR04zmoa4AFjutwTr00Ixz/KAZdW6GHvTA0zaj+cyDoAYFkIyCKJT4xJ/dhgeocT1FI2AbWOgvi/MbafzuIhBiAl1rPYff4z34cCf+AFlZrNhdfDbR/bjemD0wACzok75k+lN7Y/2nMxDiA8Q93OGwqSr88nqx9XyGHK7ngVMrGAHkgO+kfVELX6AAurMz8ewogIUEj0rRo8qeHGR5BgEk+735vQQ5PP9dycMR4gz4Re8vlyxic0ahtkua5yVKnb0F05sAgthCHcKQb0EoAQM3gC7Ao4uBLeiAukXK8cHX4N16fPcRDfhkNiwMiAtfGEhwSEOOAQGIiBejGMzWAQqUEPJg1gIRtPgFIn5RixMoYQthePnLsRCGM9AA5C/Qgb9Zp3OdUyAMGHj5vmlgDVo0QuPf9EaPA+CNDQ+UG9dQhQ70DXOYk4MGtVg21oEpciRvnQI753l0lXBdHesY44BoRCNUcfaiE/QaJwi5Ds6ghDrUYQtCoAEiToAIq+fX0hhYQRLWAWVhdMPPXfayCKixgjhPufH0qIGfjQr4JJxDzhVwxjkwj/n/OTfDGZ3//DlAv/nLZ/7ypj9HDQC/AgzkFwUvR+7PWWcDTcrIDKx7NNaVrftamFfkWx+51S8RiJ/LHLkyr/ruWZzzG9i+9q0L9MhFjoIAFKMR1Sd67nSQ7zrIPAyewIJKcy/+Mbie9sy/weyr0N/cezzEKCDyz2FPCHIogXXNNz8OwiD9q7Nf9/QcMhbAXgCGgQ5gnd4doPs5CpIt4DzVAjlokhlkku1RgA4IQQUigQUKwRaswBYMHAduQSZsgSZIgZF8EhzYQSqdksJ918KtQSqh4HbBIBxMg8KdUipdnHqpwsrRgJL1IC0ggioEoSqkQgRUoBBoghIowREKwd31/yAN9BuJDdiAUYAgIEIEIAIW/sIQqgIteJPGAQI6AMI1iOEXUtfFqQISGKEmLKESnAAtvGExgNgvKZkO1NwTDtgKUEAeSiEH6sA1GBTCYdxBDSJ1pUEqqMIBnoAOmIsUREAcaCEtZAOILcAvCMENOMEKrIBzOZngVYCUNV7jfWIFCMMoemIoguKUVdmUOUPjsaIrmh4rSoHprSIqNp4wZOIoroMrCIKSKYEgCIIm/OIWNAGJBRx0hYEb0kIcvmEtvCGI0SENLIAdnkDJ6YA7/KIgkMMvKmEtqIIkMuMWGKMxEqAi8mDNNWMjdGEXXoM16IAOKME7CkESusPdMaMy3v/jyulAOIpjdAmBKpicM8ZhMfyCDmjjL14jv70jdD2XOK6ABfJgMy4jiN0jLbzjLxqkILhDG57cD6oCJP6jHZJfHerAJdSCNygBwA0CwIVDdEVAI56AS7qkDqwhTTIhEqRhBHxSGmxXKXnXNHwXw7Wgdw1ld60gUR7l3hhJHKQCEapCBDjlEOpCKrDCVEJCuSwAIyKBFJwAVEYALSyAJmRCWI6lWI4gVi7ACaDlR6qdKlwDOJRdIfakC0oDJFglImzlVmKLKqCDN0YiyqGc3l3hTGaCIIilYSaBCJ5AQRGUTgqJY2IcHPxNKulCGkjDUsbBEMZAKsDBArADO9jAHyj/giLYQCZMXhLUQBKkppMF3iaUIim+pmsKnmy+ZidCmZSRopTlpinqJm+W4m265ijWgCtEmWymHhJAnQ4sgA6koRCMAgg+5xbUQAhqwgl4UzZ4Y18KIWDmHXdqYd5ZYBqGpzty4dChwyEKQQhugXpCp93B5AH+ghaqXRiq3XWdgH2eAF6mJVd609M9HV8ioj5G53rWgHoiASQcYhBepyRmQxFmYAUup31qYGmu5weCoH1a4RA+3XUOHRcCgiIy54Na4AkcIlOW6BbmHQ/+wgHSgipYg/+oZ4Vy4CiwAg+wgo3WKCTUWQQ0w45GQAT8wI+ywgnK5QrSoHfZw3chaQMs/ymTNqmTPikL7g0csIJU6gIrSAOVUmYq8EAEWKWPAimQlmiN+igFVYAUaKVWSgGQ+qhVHihfmqd5ggMrQKY0wMEjwME3GGV3RcOV2ugpnEIE8EAqLKV5Pl2JHugpEOGZLiqayiJMMiXZUebfDGUNGukaPILCOYMTUIstdGqn/gGo/oETOIErdANPoaZ0ouppJoETJAM7RFBq5uLgyeZqCoOTZQJioKatCgM9rEPgzSqwzqawrqavCmdq2qqv2uogiIArGGgj8qgUnClYVACyUGsjSuU1pEK2csNepgI6xIAqHOiBaiYkcENd+miXoqtVlmgqgAM4pAJYIAG13uS8Iv/BU/KAZnZpu6aCVEYqZhJhjvLAgUbAVMbBW77loL6lS94kwzZsokolN3hrKkQsOvjoS8bkCdTlmSKBMDBsx9LrDwwspGoryW6rj8JkI6asj0asleICK9gBK3BrKgxsuBLhIVYsBnKsznbsApgSDVrqI0zDIwzt0AptDdYgeLGg0hLlkjItkzrckkJtAzhceDFc1NbgnTrc0Q4tLjzCKeAC2L4D2NrBI5DtGrDCKfwAD6itP5yCP7wtLmCDy+JCjeYYlfapNOhCNGCqwuWp3+rp0ebpnaIgvxauNIDt1+JCNLRt26qt2nbpD5xCjd6tLlCmHawgknrXktoCtYSALXj/ruf+gRl0w5Rtwq6mZjesqqqiJuChajeYQTL0guz2Qj6Qgu26qg1sQq2qZhJoIjVsYuAFb7IGL7LubjdQgxmYJu/CbjKQQi+QQjI4wZitQDggAdiyQuMCKpD6QwT4w1/4g5VWaeFWKS7YgeKWr+JSKdi27df6Aw/4A42aL5aG74/+APf+gP3ibwScwss+wt5GAy5gKcZJw6BSppDy5JD8Dd/s5E5SJjdIQ9vub6DqL/7iaZAQcBzELCvgAv/6w9zCL/+6LQX/KAnj7yME8Mvq7ZXqggD3KY2mLf9iL43a6AkKrdBOaWRaqY3aaOVGw9r+qDOAKY/+wOBIQA98gSrA/4HG1QIWAI0TA80HsEKTfkMkaIgVIwQgEOU9MKk9KDE3iRKgxIHmNsCOWPExAAAgKGmTssIrvUARFMEXfIoARMISk1egBEotWAN3DeU1TMoLSMCX6NYd0EA0MKnmwoEATMIxeMEDaAEMSMAjIwqi3ME1OG0DIPIyAMEyPMAyoPGRMukWIMB+uIAHkLILLMIiYIA0MOk3MOk9cMMXKMMLAIEKAIEEfIE3ZNd2JS0cNAKPAMAUaIEEdAAqoMIRHbOHhMIGdEAHoEgBdMAzR3OK4MjPau4lqEAOZHM2CwAKekOPJERPtnIDZEKIFJEYJQACvAAmSIAV5IAWaMEDPAAQsP+ABNTzEsBAB5hCMSfAHJhAAvizCdzAKTRAUDbATzZpPUzDGSxBCSyBDDD0EmQIyHxBAKwykwpBGk3AAEyAH/gBM78AAAhASDNSF7xC0YRHeNiJFDSp1DrczzYARnPBBIAESHCBHCgBkzJcPcCBEqSEQy+BO39BI3DXFi9cA0jB6hQWjRAWBgx0A0iDN3xBEdSzDFzABMgJeZSCBojCVg9DF9yA5m6xP1AAAzDAInAAG3AAJzCAHETAkv4CCpCTQ1zABbSAWaO1KbABG2wANMiCBhzAXwe2Bnw1OUHyHcDAC6QX0uHBB8wHSMzHIrzHAFBAKjRtA+hCAIS0ZiPEULv/MhengTd4wx37WCSkQZOWsRUDQCMcdJNKgxIAcj3XMxwnBB68QByHkwCADB54wyprbhzgAQAAgS1DMgvcASIYNZP+NiMzsiMfiiTDwB3cASRYNpNiMhDI8zJgQiRs8RYbNAXwhwuENyqE96jUQSFTN3g1whcAAQwUgHsfgnuriBvQQHWDE0IAQC2rQAGgQjKLiIcoACoMQDNDMzN3wCEU+CEQgQ54V55usS9gszbnQAB8AxwoREj7CHd91zdQAD9fjD/z8xxQAB5gAgssAVC7sxaoAAzIQCRLQAFMgCksQiigQocrQB5sw0pbrUE76U7rAAschwwcxxJIAAB8QZEH/8AeN8A3hMEENLmTN3kHqABtCwAK4MArDA1Kp7QHnABLPy1Bf7kS4MdMjzlb4zR1s0IdyICaM0EZNLQFCEAcJG3U2sEWzMgT04cOJG00WAMeFIFw13MHbMCH/EZ4iEIpiEICbIGX4wJZ33Var7Uc/MKSxkBc+84TVEJdc8FZ6/UG7DU0OMBfHwBgA/Zgy4EKvMCWrLgEXAIgiDYeHEJZL4JZ50d+TAAF4MKSbnE2AIAyMPIy9DoARIIuJK2Of4M1XEJuN5FfAQIc1MMKSsPuAIoAZLEhL2k0KMFhrziiyHYca8kdvNJt4/J5dxcc0IJIA4Cf13MPIIJlM7g1fMGvy/+zCqg5i7P4JLP7d1X3JWACECjDdWOCNzDtI9yAB4z3jB88KQvCuOv4PdSCcJdAASRCxEdzIsx30qaBQiEEJmSzi9PVh2AMyH/IBBS4DORCIiSCDLDADlTDJFSDF5TDJJSDF7B8ORwDzMv8zcf8JGCCzsO8y+N8y7+8zjOyMizRCKhEiZdADgx5fMtAATj9BKByeM/4x3uAEDip1P6ks/t4Qwd5kPcAJkx0AEixd7ECIWj0k0O5bRc5ALwAA7yCCRA6Sv8GNUCCkSatd0ntFmuCdDAAB0wAB2yEgnv2w0WBDDABEzwBE7SCDPQAHtBCtdcDEuAArUf2fKzaQG/xI7z/+1QDwSybCCe4QCi4wD8TugesdN43AC5gAEekNRvoBwe09aRXupvQdSW0gOvvtaf79agL9ldLwAvIwAdkTQ+wutKBABGgsgfoxyK8/iIgAAaYdtLWAiYowwM4gjw/AAAEQCXnetI+QmaLdI9w/xg3ACgtBGd3d75LQx3AwPA/vZbIgAr4+yEQluHcAfAn9ioXNRwARLZIAQQAEPClyJc4DRg2vOetiCMgQLTkKOCmgIyMbmDAoLGmYcM1l4BMoQjEggA4DewxPHXDRShUCkIpQCXTgyaQDB81/FZLBRAWBRIV6HCoQwEiH04wXMMtAB4BAjDlsCLhAjQFWxMomMPp/5AFL16ULSvnpdyxs2vRop2U9iwmtV7kxnXLFi7auXn5ol2mrC3gcpOqlRvhpmiiCRtcuFjUuHEoD1sa1Gs4rXKDnQ0WsJBRogzoEiyKvMHzJUC0hpA+TJjA4LXrCURefPli4UsPbV14d3HgoHcXHNJC9uSpufIaQQMYNHfOgIiOkAxZRZHxhMkFJthZvKm1ucFLmqEaL1qE4EbTBvcaTKv1AogEFRIkvDYfGVUCEQlunMrM/hsMOOGAE1PYMJADOZpag4dafAkABBgqmbADDjhgg40NMoTmFQ0O+LCdA3zwwQEcXnhBI43u8MWaSwJ4QQ4XOIEsJg9cQACDneoZaf8ZICSS6AEAAlBlDZCMa4AVPIrA5AsAmhQSEJEa4GYggqYC5BspG0jjDDc+wOiDiwqQYKIOEEBggAGIIMINLF6ABLkG4AAEEFqqnEqANNhjj6GHJlJDi4qeKIDQAsL0UoeVphupiBwCrUgllhiKgJqattqqJsmEAK+hR/BQQYuhOhh1VCI6+EA6zVgBpBhvirlEhRxyYEIbP6Ioh62yztL1mLKU6bWtcsyiS62/zOr12F93nUtZZIXV9S9mh9WVrAcA87WwSQDQFpNDZmRDRhc8yHE65DY7oYfP1C2DBRB2AeCNAFYCKQICYLs3NgKKSMiCItyA5rffSvnNN/6kscz/siNb0nEL5hBojoPmCJCi3Oqe0O6CjJno4Y1L4LCMoRUS6CIBExJIgLxFMFBtvQZSQeGF+eiDgQsGzLsvppgwwAyklr7ZgoELTdkAwQHUiwBmC9Kt5IIJJxD6QMY6PCDEEH04oBQEXgik0ALu0MEbF18YgDyZzC6P3MrSwKOkk7QAAjVV4ADQKR1ekKAIvPctAg9uzF0jlTsJWqiBLBtKow4wuz4EhiWJKI8TmweQAwv1NEtDoEga8SaSztHZaeHCA/izIgkITSopIgj1hJVy16hFGTUoghSknSrw4NKudFfAg1SPAykVECTIoQSjOvCD1KSkuwcOVaIqCAAW+FDh/4EpylHG2uyxLwuIB7wfIRYVyDK2LEyixcSvtY6RS5nr/7p+fLzaqgZeAHYR4P6p8sffyv2nMsggeBJALhDggUVQgGXlCkkEesCEMjBBBg6UgQXe8IU3eENRnCHCwxhQs+YMgBBfAMEb+vWBOYjCAaIohQpR6IAEUGANe2qAwjLTAFw0QQ430GEOdUgAIRQuThbD2AX2cAEYWGAXaTDcKfohChWO4zcmQwDFLMMeSNyNPhJYQgHuYyManUcHIGEPZhogiDNZ6EAH4kKqkPYCC0RBQhOqRAs4oCEMoWIDJvBQ1T50AFF4QAIvMEoBDuGGFwhAKmfggkxo0shQhGIRW//YzDVAUBFL5gBuAaDFTowTjTN05A4woM988EAcpzRAF5EQAEECEADCnfIecbjEQZyEh0tcIxXesEAOOhCTmciEE4sYgBJa1oA4BGAgyUTm504Jkm8EABPVq4hFkJK8NXkiFcVsmSoAMJG35SBSLWmAMESggATM4WTp5B3FOtUQVVhgBDkYSgs6MIEODOCeRDhDDKNBCwG8IRCxmIL1plC9klQve9YzjCXEkYuBPqAc1rqeRCPaPl+5z6Lay96zNLo97U20e9ubaEQjWlDsmTR7csEEAFgaCD/cAE7IsYyRGvKLdEWQCRCUgQpAIEJaZIk9SJDDc5wzAE/gAQQg6Nf/IUwwjlJoQBRQdaooErCChrTkSD1B2CkIwMGImYIBnCDACYoERBt64mKtyJh2joiCV2JgHFH1kAag2AVX9ESGJ5CAKGWwBBh0gDFlyxl5cEBW5IhTB3Lwg2uaEzkEKIFeMFNBD4rXtAJUYjEbYAwe9Ug1z35IA6HogSCPkpQoWMkTCOCKORWgjq1wgjJ9eo+sZHWVTG6yTwyBBCEIFSYZyIA+pZwOK6y0SgHEgU9xAoQSYPCloqDODRKwQiU2MAfWYsoFMGRINKzxBQG2MhK64CRy7BAJAPTqARS5QPJK1QFC+Mdw7sTERCaSAwCkATnT2EI5T2Yyk3UFAZabYctO//ACFvi1ABNY7GKP5wcsRKMeaahFDwSqhoE+dArKKOiGqzeFWHQiGBieqEXLkWGPnrgab6jGSQ0zAg4XtKS4QihBR2CIYFhiBrjK8IbVYAhgGGKgGp4xRCmqrR1UIYwNAVmcXIaiB+Z0OzmwQFKtARLLaII5QdMyAuRwBjxM2QIWIIIJhqEBuh7AzE7MAwYcMuDjbNVeAzIFgcJKgJiGBBdnuFjT1tpWwkXAA2ZGM5qhCg9hMARkduhSRmQAgwRvgBMeKOAiPFBpD+AgAiEx3AlygRQ5MJYLXIBsA9qogiiUoBJ7kGMLMqRZzl7NaiJqhwYSYMhEkOoQsfiCVAjhAv/rpjMB8NjKZBpiB1q4MWY5iBUSBVCLuUmqAScgwKiQ0tsPfMRcqCzItgUAiNDtJA4vCKVGBtmB6FpkA+cEdldukAojWSMArgLENeKQhjTYYQ2YSe4jAGElACzjAcUblT1HNYAPIEKbDElFox6lBgDoIr8Y2M8rTNCFio8sATiIae0agq4SLIEPlEiECkbQA0IYAwtYwMAv4BAHJfRABReW+YXbtuMR8GGgJS6xhne+YcPwAQ3W28EIgmEINFSBChkAcvVKrIZgBKMKxtjBG57eCUNU4ehVSEEQRlBjG3u9ClUYgiRu0QdJAGMEBvX5i3FVDWMoIb40tIwdQMCCEkD/eTsSmDIIrlG7NTQMYs/xgxJqkdSkiqOpcvVBmkWx5jZntT2VgcQNwrqINFroA/7BzDSAZ4w9M41pR+R7kSjQBUHPFarU8E+c6jWqcm/AkZfKFAEOdliGnIC3p6unH/ygA8yUOgo9uCwlKkH8OroaGia4Wh/7qIE8EOIFRLAn8grQ0y/IAZ3r/m8o2KzwumtxCUuQJwUFQAtFsWcNQpDD8epZqoMnlyHgKO5UGpHBw4Fg3F0z9/Coa4I5/DedQkETbo+3OoI+gKAIACAbtGRLAEFzWmkqLIAFMGJU6GkADsF3cksVhEcFgkIFvkAVLoMCTsbieuPicCCb2kkzxoAF/8qgDGQgEbhgArSBFwRqBNQgB9TgBlVADUqgFVyMB2MuBy7Mwi7s5mTuAYwh7MIO6tCACpzQCVOgEMBAESTBCqmg6KAQ656QC9EAGCRBEQphCq9gCLiQCs7wDMeuCW4hBPqgDUPgFiSBClysxqjAEjIgCKhgBkbgoKag68hiBwIhEEbgGcghFbKkJezgU4jngcrgCVjgBUAABfyGIXCBAmqGAxaBCzjhYaLjPSzgRDhBFOLKzBYPqmiNMuxhDVqCjCIPM+oBEuRgEy/E8giEEHqiJ3aCFchhrVIt9FTgBaoMCRKgzOaK0LrAqhjCZ8IAAWTDnhgg+3anKxTABbrvqv80A/cwotwOITowAxfC5hJ8AQSeIBeIb0JaYGhcABWSb/mYb9a6gBCioJ5c4yhw4/pKpuJeoQRP5gpGoSFSwcCW4MAG0l1sSVESURD84NMWDJ8+4M7c6d+0haUiAb9CYg3iAAX2CgbcgNwSAbhyoP8qTiRJRgFiSwo+oANujVBEqQi+AzPESU4AwRo2p0qUhD5OBymIYNSYTBVe4OPKIAeWwAJoQVJwwRVI0ASAozcM5pTEyZNKQAYeCLOeJjZk0A+UMBZmQA1Ibghy4QZ1MBhGIOaKcAosTAnbsOwkgRSggC3b0i2hIB/yIQ/yoRd6gR3YQRHesA/2Ei3dsBv6YAH/xqAb3vAPFEERwAAMppAdruAuGYEdnMAJ2IEKJWEIyMAKDeAM0SAIbGygRiAXDMEAGEocyAE8egY5foIiZCX8ZIAFkAgF0IFPuCqsMpFALIQAIqDwQFECOKEYFw/NTFEE9MAp0K/NyCgCboALIiZy5owBwuBIGoIVwqBpJoTPjugFaIEVbkDQQITQ2m066oUN6AysFCApTQAegM2cEOCHiLMl6gH3CiUpDoFQsO2YmkSp+GA6z3EWoGEDoAEaEqAUmK/5XuED5HECWkDBwuINisAPTIDiAsY3eEMAO+7USgAG7G40kMiWQCc8MEDBZGMAFOwDCGczaGG+rGUZhMQO/6ZjGuJAeDritwrgAhjnBbRABhjAZHjDAfTxZHaGMwjgQztADlTnDjJtM0BCFxqhc5AJAg8ib/ZKBuRzn4qjyT5jNEpABYgSM/zhBpCyN3iUAqREF63DgZggwV6jZmJj8HTBF6qAF3JhD3MBB8agCoqOCvLQEgxhBHYgB7eSEGhAF3SBB3CBFViBB8ABHH5hCyjABhi1EK7gD7qhG1ZgAR4BF3hAUHUBF+wAUwd1UFnhUg0VFzZVF0IACq6ACsbuGYYAChjBGdYgBsLBBrohBnhgDOQQDdHACfPQAFIAMw0gD8WODJogBVsidH5CGRwBUKxiCVRgB/BgF17pOAkEQf/CcxE+IBWOzQIkoAegoRgHTQNmzQdCQTqWLCTGiCGkYABm4TnYgAEQ4BlacSdwQTpBjzrD5wUuYRQSYNA+5Gp8QARSJbm2AAHSaGg2IB2cqBQGphQc9GRgqmXYwzgiIEzkMz7nE0m94X+iRwYyJtUogdX6s7qGQUBB6xXiEQYbLCx2oAhw4BV+QxYCphR4wwN+6PZaECpdcDSm7gs8RhnX4BHgQBrsLQ2kAQ7gYA3gIBpyETl+IVa0YAokIlKcKSZfFAZiNEWCYgkmoGR01AFKAR66gAIwQ/2ckQvShBAQDtEaot9ayW3ddpZ2AQ/eAATOIAqUwJQYIkvs4AWe4AX/oZIFfKEhmsFlR6Y891G7bK8BEMEYcKoVEmwWwKqDYGMCNiUbAsENYsEKbvAGjYEKDCALSKAQhgAYDMAASPfHQgzq+kAwW3cMBHMBYkBQL5V2QdVTafd2WYFTL1VQOVVQDXV2CzUwu2EMWPd1WbcP/qAMzxAzgSEFsuDHuo4X4iGqnEgEBvA4srdwaGEHHiVQMMkgnI1PpAAHGIANOMGOCCQMokEXlErcFMDMjNEHxJVcWSLfIo8heCZdyzfwOogLPGFe4gQXeJFpKEHVLiB8ogAEEIBkQ4Q7ReEGYigkXsLyWq0momrWpOo3EiAPKOAdpMQ4dkspjKLaMBAzUqlJ/y1gCVwwp1Qt1DiBDUKhC0oWzeAxEITC0QgFN4oAAV42hVZohX7DA9gJDs4ggu6uEVuzp3yBZSxjOd51cicAAfzgDBjQ4wRSVu5LStKgEcQNBnoABu5AjAnBkI7BAgoAnXwDQrugPxoAy/CFct9LS9bAGrhtKiDwvDABE/YFGF+gIkPCDlAAO3LqEWlAUpDAAwKGYEpQAawxe0/ADbaDCfYgwRgArCKmObhAECQMBHrAKzl3Bu7UAEo3CIDVlEs5CCShEChAUHmABwxVVF/5dmcZd2tZlkPVU2eXlncZF3QhAkLAHcbgF2JAlT83CI55DkdgBrRBFqDqGJPRzSRlJ/9ooQdkRQsARXaEpBiejTNwAGpMQUYYoA7ggBVQABTdYA7id9BCRAPGFbIQBn8jbyfMyHzpzH/rQDX8zobI4bL2wBwrIYEJ4RVgrfkOIBQohj2qiHzBxQVcbQ58AB/6iJ01ADh8tJlcghBurb2U4gVUIw3u5CBITiDvjgkqRLPmwAFouB1s+BiKAAhyQALuwCC+oIdjdqpKAYpEgRqagSGkIQoGWTsgiAV2YIkTaBowIMvAyhRqJjqY7PYaCCpHYxcgTiSc5wVgIBZSJCMK4IiUwUbzw2sHRhZwwB8aIAyyjKjkOLfkBA+WwQsk0iCK4SCUAQjoughYFg/+2CdoAAb/SoAPtkMGUGAnkkABWAinByYpe0dRqoglaCAQJotbWaAFgiYTLbk5wiAVLsECAkEcflAFbswAis500eDpSneUTZmUT/sIrmAMXtkfChWWZTmWCRWXY9tQOfW2e7lTY1uXRdUOFuAKrkASUPmUk1kNKGEVwJXQSuEGrpFTGkAVKOvjxM9RoAR0hGAANhGcweU8IEsX7CYKPkD5aNjMoMETCIcVXTEktgCGXSBDMIQDRI3jxGmAp/Of+WCvOKFfm28ctGvJ9KtANIs/UcEEPquPTLELNGHJTNMecEEKEOEEEEEHLkEHIBwScMGYqqSVvuClrSD8Pq4EKoQDko+GfWAc/zAABZxkffYlAADhEnBgZH74FFcI0xiCB8jhDoyBBWIBq79YqUCABl7JEonKORzSiu8AO4L6BahaM+CAFl4EI7RaI7raCkqADUZGjcV6iNcAAzgorVOwmKThBZTNER7AC45BSDQbJeirX74gDb6NISZsCUrg7mTgBRSlBoixetPsN0JBEJ77HgR5zwjlacLT0MPqAyJgF3og15R5BsJyBtDAdE13CEy3dC99lIEB00s5tZ23EBThD5yADLrBlTNVtk/d1FtZljN1AcLhCgrhV4mb008ZWC3hB3WQEuiAZI0xfj1g9TjuOVPBE5jgr9mlBHIAE1yprOxBCRYLYoRmAP/C6LtP5AOmho/Y+QA4wQ2+AzmSC/7YG301qz/ZAAGSLHtZwRgsS44q4QkkgAhegfmIwV9F4AcsMjwoQEMGHBrmAN5Llp0TAAlC4hV1a9pGBXmQpwPOgDjSgE4aARAagSSYNSib1ROymxMSwDe5k64ogAa84W0vwRrg4BpgwpwGxoniahgQIAowYRfGUWPWSgZ64MeX2JVOgPLmzF0jR5xb55Q0YwE87wmegA+eoAcQjvMe4RqmQvjks1AwAgZAABMqggHwkTcGxgEUQBN+YAsIQT67nhDCQAjqfW0X1xgslAVGIFCUwUnkg+3jAwhe4BoGXowA4QswIcyiIApegHD/Sk8U4kEBeMESeIEOqDcUNiW5WkIXBBnKmmYWLqQ2I2cbuGAf+GAPS0CZldkSfLXSN98AJAEJHuEbcOERTuEH9EAP6OH0Ux/1UX8FzMAGQsAWYL8JYp/2Zb/2bx8MzIAe6EEYVl/16aEGXGEbTHvSi990LSHERsAKKAEaMt6z2FkE1AOe1/oUnmGttOMzVCAAmEkzEnIeOwisFEQzaOAFeoAIHICgHZjQwAIF7E+BHkFAWk3cOVHAjIMVrN9j5YjoPaAdAeKAwAMOKDQ4uKZBvQZIhmzYAA3iBgUODvgYeHGgiAgJEyI8CImAnwF+WpTs4OcMrUgBAgh4KQAAkCVW/3JYoZlDRaIJXBT40ADU4gENBxAEOgbgWBGkAaKdIsBlkQsFCbp0EeWg1KJAyqaMuHBhD1iwJSRYUGHBwps3mHbA4MLAFAc2HDhxYABjRxFfaQ4ePOEGLKWwTFTgqXUJxBsQX2B0eNyhQKICBdyAwKRFy4Q58ExYLeXAQYIVJ24wuEvXLgNCpxp4PEjDzZMLTJiUKZGjmgU3MmQsWSIh+AtvHRvYa/AN0JcHjhzlyGEhToNprkRsy0WJEq/sufYhWNDgnt+DrEDAKGG71YUJc02xYaONF58ZsWaUsM/HQIr9/PsbGNKEMMIkIQw99CRRgytmUGPGCv488siD71SABP8PP/AQQwjs/GFLE7aE0GGIINrCDhjhIPHOhN2Eo6ArrtRATw1miGMAMAbcaOONOgIzwwhWjNCJNnMEJVA7GHUhxEELvfYNeeRcMBgllrRwQQ94pOJaA6cIQgEGFHzwASEUEBIGJK6d8MILRIhClJEDDaUBJ5W80FdCj4zn1yMYcMLGQ36ygcMJ44nXACvkzBZWonwkIktGGB2gAHgHHXfQCpxsoE1E0EBjwkVuvjmUBy/QkAahWTYAyQ0TrMoqSncA4NJLsQKgBU1L5HDrEsrA0AIDcwxTigZsavBTnFEcswxSSjWVihIvOFtHHZ5gAeYHd7wBgAUs5HIBt5WQFYX/BS9YEMgO5qpQAAMMsOHeInRxwcJaO7TVVhE9PCHWYJXIoEIROywGQlpu8LSqH5A9oYIymbUwRwIJmGCCA569gkAPfsTFgF2qEXINnvcANtZYJajwAmSUwQCDBD1cAodfCdUTBwCTHOPFAw98IV0DNySwjyWWaJdd0JTkIs4ASqxxzxq/RCFDCWU8zUQis+yTSywltDID1q10sk8GGQyRQQpGkODEGAvEcPYCEUQQA9s/tO1PBDzIHUEFwqT4yDsQ+rOJMzzMjSGGmzjhxAJ/Bx5D4IfPvckm7+DySDOZSHGK3IlbjmEMmq9wxRVVBDPCCHwww+krXYiQgAjwoC6C/zoYDBreQXZgUEUPI/Q4gxWtUBLLLlgeFAEBE/gxfPF+fPA7IihEgcAwRD0/EFAMJNLD7w3cief1e/bp5wZs3GBmlpTi8qS3iSYyh1ACASWKKDhAssY08cPhSxRcsBERKhuggkqnoL45jAGY6w0W2IFa1LIDFfRKXQzgSQsmAIMvwGSCMhnBb3JgwREoQycTQEVo2icsYYmCCypYBhCWUQQUCgAOEbjBAHAwgEUgYBFSmQoBACCAL7AAURf4VgFYEAUVBIJc5sKExeiCxLlwgAs9+Ne8nIgJ0X1LX4UxoAHFhS72qKtgLUgECx5gBS0wzGFd8IxVusCJOzzQFKfhgP9cGBALC1TDGPvYBy+4wItZMGMVLdAXDF4ggTuojGRF2IU3rhGHO4lHftGIAx684IVJlMMLAJAOLnbGCGRochUQuAIvfPazoO2BEnt4AiXsmAte8IIF92klHyyRgSxkoBCxnCUJbLCACixAbWqTmzMi8Mteti0Gb3NG2xaQiR9ADhsQesQPNCEFwF0OcHLjATgS9ze6URNw/ljACiLQzEckIQnaZFsMIME2uo3hCoUABh9ysQofXMRRQLmBLmggDkKErgS36yfuRhALXrRgD7FAASuyJAU5cGECDZzAAIYXhmjUYw2pEMALuBAUI31KWFyoBAwEdRBFKsQvuKAAJzj/ERHvuYANckDERwhlqFxMUaYXYIAshjIQI2lAAXdQgRXLFQhKLJQLXOBAXdiQDqL8z0gJOMQUzAUCc+2gXAm8X2q2yAU3SBCHFAQCC5ZQArAuYQRAwAQmilCALjhAFKVoH1bcpxcgFGGuRRBAGkozAATEMIYzZMAiPFGMSOBBBSVADxPGIoEgDjEQUd1BLPzArsi6hw1+QItUC1jAe00RSkzIgVQXqwJCcEFjbuSJH2IBhBxooRLQcFhnyljGNBKPgXFZIgsKaC5x7GMbq6DDKpDhNV7YcbjCFS4ztMEFP9xhF5HIBiCciw5ACACSkqRkAADhCxwo4BW+RUYb2gCB//CK97cQEAMzUsAMXuSCD61o7wyCYYmueU2WstxGFuSRhSwgIw8hMNsu/xsBXgZ4wGmLwSicoIgQhKMCj8MGLhzsD1wgQRjljNs2EzdNbU7zcv5o2wqcgQtcRNgZmUiChpqguXSibRPsKMQQUjCETgRjBrwwxAzsc2Mc36dHhogv2IawDX5QbWhPQIEu/IIEHLTxNET1Qx08koYAvAABshiGD4aRDi7kgsZzSIcfKvEEJeRpzPWYhj9OAQlEnAAREYAEJFKhi2jcaRojbQD5ClCJSiQizx0wAfSep4EuEAEITz3XDo7IvfyhohT/Wx+kjGFFn2L2XBN4T5/cY9RDFP8BAF8AAA4/XYSvhnXUWgCACjrABlmsta1tXSsO3lCEFwDBArHGQxx0AEMZypABM0QADpQQhzgE4BhT0AKuyiCDWKggXEMMl7meMNpFeC+ysziEFSed2Sd8qxJ7qAQTylVA0B4iYxkzqrq4UIAcwGAJF4BGF6oC7zK6wA0deCBDtdgCn7aFgAbkRTpAkQdQ9AIUdCA4wA+eBxKQAAKrkEfPQBe6EXhlCmqguMXVgHE1hO7G7c3Odj5uie308eMZOEIhjoDy/NaSvrNUeSGy8HI6gGETC/Dvf3npDAEHM8AhSIYN/FbzEITABooAAxhIwQ52fGLpnzACGIwAdSN8ghT/Ua86KZZOCqpbvelVl3rU2dENthV4AU1gxBCMALYUeM0AsZixAerotVrGvRCepESeC2D3C6DADn4ZxWjrYlTTKuEXGCBEE1WgcTW81xKtyAU0hiGKV3y5AFHoi0LggIhaHPQgCX3PBlzgvQ2YggiqWAMuaLALzFpA25XIRQsqQYlZOA+nxGKTBxJWwKgWMBZcCL2fUKGAYSwVThX76bXN1QOiKt+0E+hADwCALTxwOiahFuuoVVANALiBAa9YNVtFcRUEgAAIEgCCrCVga1xPQNe95vUAdJAGYcfE08cAggpUgAkLBGz/BRy3XdjAJ6bACVnlL5dlRSOgbT3UQ08w/wI/RS6hZVWWhmmJUAJPUAasJTGwBW+hUACP4VCswgUdoBaYsBYFpAKxMDTY0VsBx4KgkA8HN3CgoHAQ0AYm5zUwph//oSMpoCND8B9qlwH41QbIEF4LZ4QQcIQ0CAHedQRiAHMqx3L0lV9ZcARUSAeFYzZIsEtSAGALkHMEhjYRsAKMYANj4AzY4GAQhg3+8A5s+CARBmG48A52sAJPV3XOACHY8A2bAAZcBwYhsIZtGCFr6A8/0A2ZEGALEA5mEA7/5QSMYARxJ0vzFTbB0ArvJA5VgAJjEAjk4HoCJVwtYEfi8DPtxQfBwAdocIrwZQBhEzY8CIv6YQi8sAqQJ/8Kw5AAk5cLKqAY4DZVVsR7SNQnlsYLaWF8Z8F6eFYJDPMTtNcOgUYIylANT8RvuTAL77FSDwENQ9Im0TMUoiAHknZ8khYIkBVZ7zEXftAD+bcDivEGXwBrLMBKYFVYOYAJACABExAxoDEOpVAKasUJFiABKSMBKiABX3ANQoADvcZ+MnQDKBB/LuFpMkORsbILBERAFuB/gJca6nh8k3YvufAE3FIAfNBE+jdE4yJa/yeAAsgAh1AC27YBsqBWVrGBj0EEBjMAHTA8ibAD2ccWawFQ+tJDBXABMNADgcAJ80AHeVBwBRdwvTCDJKBJMDcEL+aDPJiVOqiVMDYE+SX/BmJQhEg4lUgoXjTYBmJQg1VIS1E4hVVoXyiXDGRgc0KwSznHhTm3S2C4ACHgBJvAAyIWiG8oYhFSmBGmNw/CTI8TYW4YIRHShm0omP5AmZR5CptgA92ANpnQDTe3AJswBuGQB6SQX18ZS1T4llkQl/JQhWKQciiHcvwAmzXommnpmkcgD/ZlX/SFla/wCm+1VrLAgUbJgNiWQMD4dy4QgHRxCERkggakAvjiLbmQakEBaKKwDWpRDW+wnW1hAbywLu7BCdnIjdYJJ9Aojr4IbirgB+2xUkjkkWnxAvsHAqFWWIUlVpsGAAUQMaExDlkBkBYgAHjQEiwRCdagBAuJ/wC9tqALegOXEGwBMJETKgCNYA0sESsEdDGLQG6cgACccAiBsBgDhFlvEAWx8ATaVgC5IAMnCQKMNUSEMACcUG4cSqOHwALbZgqh4QBXYZMJgAAdkAgdQAREajBEYAGfBn2YoAIyABbcwi1VEggvcAjRdlKcoA2vwJQIN4NLyJZph5UwJqZhmgVfSYVqCV5meYRJCF7fFZYpR0svJ0tySoWsqV95YANIoIVa6Jl36YUCpjZmYAM/UIiUCZlueJiJSphvSJlt2KiVCan+kARmoJl/enOJqEu7RHNmYwN5gAz3Vaco55quiQxvWoOn+l3e5V1oOoStqqrIcASwugrbQP8ACvCPPFqTXfAKHvAEtVGcb/AvJShVsTCj6+Iui3CjBghuFsAH3dJDHTAHwwIUIpQAhLCdwEqC0BcFfvCh5AaAnDAk0goU4yAsCtBE7YiR/6IYBtSeLNmRPVAEiwUC4zIurMQEJcAH+LkDntYDodB9XfCftxoKPUAARHAyf4QCdQBDesWwLzQABIAIaXANL/FpMSEAkZAGuhAHgAAILCEAIEAEDAUX54YAH6AW68pvahEIMJCiIvkEMlAuIPCiMyujCDCyvMYAXICjRpkLXKBW/GiTr7AIcpAIRHAIBtsBh0AIXEWxpsayKTqSTxALUcBYMqouNrpFhDBAwWoMqyD/g5qUcryZBWOqdilQpl+TXyj3XWO5pmoaXqm6lmH7hGn7lqxZCL1QhgvAp3rbpzn3hWeTBEn3BzZwBSLwAeZgDuowDuMgAskwDuyQCX3zA2tIuZX5YAvQD43rBCIAds6wczjHS/81BkhAOOEAmkgAmt1wBXmQBa4pm7V5BGnZqmqpqkrYpjS4cGcZXnQwBIGwCyL6jh8QCj36j2dkkwhQAk3zBBKALWvhvMD6BrGwQBzKQFk1ooqBvRaAooLBBd03Du1TCv/pAL3rvO4IfbzHUAiQs+qCAArwfeHbPmvlAAOrrotRvsBqAVDBazSqLtvAC00EozNbr3zABzLwBCjD/wIq8BIgwAkTYxUOYDoKQAhEIAdEQAQfUAB3AAJhAEMdPAAfPAA3ALFpIF0T9BKREAdwkAYrHH8biwIfcLRE8MFc8MGWAY9rcZE4rC0v6wYoCgNRsBgoILMy6wkKlVcDsFB6lQv3kqJ+UBXG+25dEAoDYMGHcAgw/AGe0BJb/BIW0AOxAAOxYMCxEEeMdQdyoFc0bLM0nAuKsQvuuAs9gMAJjH8CQAgewAmh4AGhsAp5sAqz2pZfaZoop0lsO5VlmbvhpZZw+oRViF9VCJswBwpXMAZmQ3N72rc3ZwMigLjq0AVO0AR9EIZqY0xnU8rAhDYxcMppQ2B/26d8q4U0t/8JrmADm6CnoLkJQrAC7MAIhZCWpeqq37W2txteyOC1vuUBC8kF22CzedWcz7sLuaAAD2y8DqMAAyCPEpDAbyAA3LwL3ZzDxuAHRJWzCDABekUIOfwGF3mRIICiTTzNXfCP4Ad+CmAMzsvO2BIIVZpXOKDGeZUAPUrNAv0K2xAFIPDG+azOIJALeXXOXMCwRADEMstYZzDEPSADBfyysXAHURATIIAADhNv1kwAclDBREAABEAIZ+AJGIAFGFAHWBAtgjDTkBCRLoHTFZrC0bAGcAAHdgAHcUADnuAJhEAIKW3BchAFu4AHCM3U67wLb/zFd+AGMOAGSbkLKCDEW+3/CQQwAHIAwh/sB0vcw25wCKsw0u+WAAqAAFV8xbngBsMRAJHgDRj6BirAAj0gj7GQ1zK7PASgVyAM1nJAAG68zuscBXfA13x9W29ACNvAxydXCC8Xp7XUli2ntmlqhAp3yEn4trL7mo0MqrfZhFmQB1fQB2Mgy7D8yk5wAMQA2/DgIiIwDj63AjSXyqwMqAH2t1yYiJa6S1qoS5hsy8WNuqq9CaMgBKOQCVdAlc79x9swBMEgojswAj2s0bFw1QhtoiMxwx8M1oSA0E6NAjegAOctAucdCgoQCqGgDerIAtqsAt8sABaJB1E9wX4gB/pNEgOQT4px3wn9xp5Axtt3/9577AHJjAOE/QKHndWL8bsyuxjw+AVvLAdz0AV50AXwcEZVIQIDcNBRLeDwmMOEANZHPMMS/QVDvNUgsDxWHcZh3NEAcJHaJdIOozqhgNIijNIEkMUEoOA3gAM3IMIE0CU2DQhbXKDXlQZrwNNrMD/cUAvzmSZ3UNRGjQeXEABMvQu+0OVdDgJRYAw9MOYdHQh4gAJZrdUooARandVNDedCbAx3YAwf4AEKkN55HgoiEAo4UNIpDSaEoAOREAmNYOiEvgs7MC6BsGxUuws0QANn8AE3QMFycAMmjdIIfd+bHghk7unGQC5AjgAeMOoLiQMwRAFz7QthIA6FsA1XsP8NtGRymV2EnM3Zbpu7RPhdsRvaLwfJrAmbhQAB/GXLlqynfBvcyL6XnpmXfxoDQhACZuAE/bACNVAD1V7tLsIg/cAgNmAD4RAOIbACmaDco9A4x53LjZPL5j4KmpAJfSACeSDMREjvxuxb21AFsUDmdM5Y930G4mDSlo7p4uAJKFDhm04Ae04VIpDnB04APdADL9ADvKjkAXAJAnDxz0DB4nDpJi3CUbDpXB7giR0Lh7Dea706ay0CHuAJaH7fl8DlKFAFAC/wHk8E7ZveKI86VOEBD3/mIg/0eIAFGx/wJk0AII8CNJD0S48Hna7vHK3vPSDiN7DnCs/nK38DH+D/42MyJnUA2Kcu5EROAQSAAYLADWnADdF1DRy7sWnQMlAO5fLDDd5wCXiQ5TqAAi+gA4NO6MUQAL6w5b4A+DTwAlQbBYdv0S8P6ainBEet9YDu41gQ5ofvCTiQ4Jef4P3gATcw9mOPAVk86IZuDYCADo1g9+vs4vOJApfgC5cw1Clt5LDfJSjQ+rvA+olR+FHwDIf/AmcA5JZ/6mAvwuRQC4AQB+AQBxqLDpEAEzh9Cd5g8WEgJo/v4wRwBkv/6Pcd6S9QBxRwAy5S7XraDFLQDBVwDuavBxWg/tWxAqjr/qu9CZmgIJzbD65Q7bAACyuA//m//wABS6DAGrAKFhwo/3AQrIUNYbnCgQEFimcELFok4kGjBxEeQnHUiGXXJV+XRpYciQdFlCieWrYMBMLXrjoXbVoMtEuAr527CGzs+LGfRgQfWL4IZAFEgACRmjJlGuUDgUMYLRI6g2ekzl1a8bB8Jk7jx44bKXD1xXNXgF0obBIhAJcAoRsegdr1MABLlEBaTZJki8cXnmdVCFC4WeXMJRqNdzWmcQlFIJY9LLP8MvjnRs44CITBgAVDGCxh6mAgc+MGhdUUMLhGEidOGtm143CDs6bBvQa9e8MBVKyRtUjenNZSlUZanGuAGjUqVuxSLV8ozljHjoJ6rROIaNRacJoQhvGisdSx/kKJEv/WOG7ggI/DjOryoc/7ikSrESD+wZ0GqCWAkmqxhpZaEBECC/NCCy2MyIpJy5cAaJgIBSVQAMFCCtzjUDUCVlPiGtl0iUOXNJyLJMUUG4kEkDgAEUKJOuoIgzTSlOiuu+/SYm+FddapQJgKKjinAj1WGCTJJF0ZxBVq+nGlH2qoQVJJKx1aaAVYVqBHmGacaeacZpr5QUxnyvwSTTDBFNPIgpR0koI6aPBFB/IoIMS19+BzIr74CInMl+0ELckXGs4I5IwXFL0uUCWqGC/PPBVEgdBLLt0QPg9wQACHTd0jB4TrLkSBKRUjYTGAM0gzj5A8wyiV0EF9OWPVunDo81P/93SQVUJCUcBCUjzxPO+9TTs9Fj4KFEWBpEGpI+mSM4QVFgslov0usmzTq5XRSi/BAldPx6XGMyEEUQJddJXYwjV3McBgi3h1UC4OadJIAw59o1lDN9166xcO2myrTRc4ooHDRNn4s6ZAGnSgQYiHaTjhQFUiUAURVU4QYgtBwhCkDkHIQZfCh1EIgwKVV3OFNdfq2GLGkXGsRT/+9MO5Ef2KAURE2bg5YT1BRpZZkO9qqaUYpBuDWAcUIFYCg9WmpqBl13S4hpsSS0yDxP74e3G2OE4g+4QFdBAiRiFOUOUXRBChrjoaeqQniXWS6JKeJFcYssgh/wY8cMCLPOcc/2cqOLwZxNt0hnHEHz88csiJfHydQTLRIxNXdKgFBXLq+Ny016gmPYyKk/6lGFqKSb2WSxZ4GgUhYv/uEh1iBrlGkJWAe9BL2p3aleBvwODCphtLej/ohrNmgXRlPGPoLZSgQXWko1MaPJRZU0144SkQpGbxkzbw4dxhDsPj9Vb2XrWp63BaO+whhBDpWmTUPX9BOK/4F1r8RwQtGjMGC6GAgGMQVC0EwRrhde8G4WjCCXRwAimYTYJCyIQmMphBQWhCE0KQwm1okwZ+9WsaDfAXChtgDxSuITe54dc01iBD3dBwDfeSTSoydjFERAARv1CFKlKRCl0MMQJSEALadP+ABCXqABEn+AUUOxYvKsprC1vQwQeTmMQTFMgaqriGKgABxlTIZmD5ssMa0sAKsukAiUtEGxCzQQs6/o9iFCMbDRaQiSuuwIp+9JgUriEiEs1GYV0zo4nwlYpr6NCHPiSbKuIwRHD4ggwiAMMfzGCGFSQhE0lIgjBCKSQhCY6UQUKlkIC0ygoAaUiuFFwsYRnLwK1gBcLQgzCQ4MfupC1tSsAgvDCwgmEWEwPuOAE6VDHHOjbzBHgsG8VogQgduENtwEzbAug4xzkiwh3CJGY4h7m/PD7zBLQQYzb6Yw1ASFAHTVQiLby4TFowU4LyEmc4BYGxOqqijtmQoCCuqTb/tMHLNcQ8KLwm+ER0ZoOe3KTjAmL0vA8K9JzoFCIkUgEJf0bxjuYMoDeE8BqSvmsLp4gAD34AiQiwNAJIkIIUnLEAKSxgplKIAb5I6MJ+qVA3LEwhwHzzL98UFWD9WgPCTDREIQqRFdFghS5YIY1UROAER8TqVU+w0VTEIBUSRAISdCkEsYYVq1LA6i+UqcxGgiMV3DCRwQyWGxuyghU8QGkEmmFVjq41iEEE4i8goVEpIEETYhWCLoUhhMOeoJFmjAMccHGwgyFVhgjDLBykoa9MsMMGtrDFH/6giNFusgZI6mQNPJmEboASlMIQxjpUmcpUyta2scWtbHN5W9kG/6m3uK3AJn4bpN3mFkk1sK3dkmDLJ1LQuRL9oCY2EV0PImGrqlBmEJWpw1QEEGMtxZhGIWHBCi7AuWzDbnpVwVgPtlcY7UUrSy8GCSBKEh1hbCQgIrDfHu53vBqdZBzui10dQkIKHsygB5PgwQgQsanaXaZVaRpTmpr3iNJtrwY1sWAh7PdiQ5wkOhgpREaSrcIxrSlauTHEMhJxxG3bGC2+G8RrcGyDGs6gEKaBi2g8osdweAQr/HEKvA7ZyLhgRRrS+FOfqhCoKjRqlH3zCKMyuTePQCor4sAKyQIZDqw4xZB/cIoxj5kHdmUFLuxAZjK1+Qd7jUCYiUxmSrq4iP+60IU0Jpubb8xwDSysRwPqgVSlSsOuLnarW1mRCjSneb/7lcKb33zEH/CgiAE22JIbQGXd9PkbDRgDGBQRAtCW2hbhsIETwvHJGmSi1SvoxqtjnYQadGMFTkhGL3pBCl07wdetvVtyRXk3UGZiSq5Q7WtDqdxhL/tuooR2KJMtDFd/stib+AM7VG0OariiAv7ggVd/oNcjNkMK5jb3fi/N4iK6tYiLviu8ecDiOI8ZvCxtdyrcmgqbntvfzkBxStE8b0a3OMBvhcQpFH7mMxPRRPeKaxGlMe5/y5SmzZCGHeygZRdPsqouBe+4NxoBmlZACiaPKeLifIohrvvgIB7/bMgjEIMIVFriuuhxNPLs4lTMe94aJWIEbmpym8LUGRJAeg++MBv9XIIuRLjBh6D+ocNAIoXfiAQABKB1ATAFEEGF8hpQ5JT/BCAOuuENILYOAABMAgBfj3IaQACEFxThC2zveiN0ofYAdL3reLjEF7wRDRXe4xovUAHS7yABGFgGEYQPtL/SIIBJeGESylABCxjPAhgwHgYvuEYK/wUHARxjGct4wAPezhve9GYLCFjEIlwge9ovAgPS2M1QdxOHLwABBhcowBMK8IECuOEDnkCECoHT961rQQsS6AAqUBGKUCgAFQqgPio2IIcOFKD73/d+AYgwfEgM+oS9oYUF/ySQA/bnIAB2gAPzmR8JOPRZN+9wxsdC8wEMfMA8dc8BLcgBR3CE1AMCpEPAJeiADQgFVEiAB0wAE3jAGzgFKSuqepgGHViCEtjAJYCBJVABALg7AAgAVsi9NVgA7puAAZgAP5iADuiAF8ADAaDBXZCDPDABB+gCB3CAUuDBLhABJOgNFroy36ChBhACcZiACWAAJpwALpADJfCNQKsHOHgBFpCBJVgCKxhAAGgEOMg9FjohKcAAqyCAD+C/LYCE3kiDSOg9CWCBAiiACZgDHhSFUtAAUdCAUhAFB7iBaTihE/IHCmAABlgEDjAFBuAEBpCDE+gNSEABC7AAFmCCC/+4gBbgAA5YBE7gADZgAxeABlnQgFE8AA0oRQ14BSKgOwnogRe4gxdQBeCADiwYgFq0xVv8gFQoKl0IAAA4BryjQbgLNKOCA+JIkadoijRAuwZQO7bzxbfTjWHsDWl4gReQACAAgtPTukiwBm+4BG8IAG8wjnAMALjrjWmIg26ECmvQGq05PyibvMrzggdQgRLwPBjAxzuIgtDTvQaAAzxAvYD0wqBaAwxAAA+QPRdQyNlbBCzAhX7sjWvovRKQgYp0AxgghDsgBE9wxN9oBL8DACB4vuiDBuwzSQWwPlTwA/D7vkMAvw9IvsJrgFpIvPbLAQFII2vou538whSqhy3/qD4IfMA5SIABAAFMyAEudL4HwEbNWwIE7ABTkL45IEqhxIE1DLR3fEcM1MASYIEy6MAQHMES9A17kILzUBAFIQ9CCEEaFIAvGAATyMEd7MEfFAEpiDIqO0ffEAI54AImLMQnjEKjsodoUAJ8LAEOHIEpAIBIsIPc+7TeQAIC6AAiGIAOGAAikAM5uL3eiAY3LAJrhAEZmABU6AK6zMM8FIUuoIB/OaFTIERDREQOWEQ5SL41UIVInEQZsMQWUETaNIUN+ERocIBRNMXj1AAHkANJjJ0XQAFJMg6nQwAWHIBFoE4cGAAK0EUV4kVnBMZGqKEqSwNwfIr/iIQ0EKpm/2Q7t2uE3ojM3mCFaly8F8DGItC6AAg8PLi7GeTPSMA9tLsGPDgGC7BGxrsDT7gEMDSqNBBQL5jHerxHzjtQa5BG3yC9gEw9L3xPFDJID1jIUFDIRfCAMFDQKMuGIgCCEhA+OWTRAriDjmwAO4gEkMRG6JM+6kPJHJ2+ywy/lmzJAqCB3mC9BvAFFbDJm/yG+NvJrvs63qghCkDJB5RAEyBKAsADTBiBHNhCK3A+38NHCXjKOVTIoLRKvNxLIfWNe4gGFNjAr9zAEsgBEcQDEnxMgAmDAXBB6mzBDlCBL9g6AQCBuEyA09RBHtRBDzDTotJLQfMNJfDLAWAALmhCRv9UAqLqjVQ4gzuIBYpcAhbIgSIwuzUYUioTBDkYAFOtRcwkAkH4swaIhkb4AhQ9QBtVgEF1gD68Q1FIAAywVFaITVOYzdpEhEGDhC94AQvoARmohAvogAkAVk4ITjbYgFA8zlIsRR9QTgLdvM+rhTgoBm/8AASYgOlkAARggAGYTu0UKl0oBqZYOxr8wtxD03pIA6ggO6awBgUdNPV8RvCU12m0xsXrvGu0TzzAg2N9gS/YTwHAA2/APd9Ig0sAgCIoAsXrgTtAhBMKtMjkvYAEgnrEQnzsgXxUBaEaPYAEAqZ8gCKIBCe9MgpIyDFdSA+oA8JrvRP0BhQtgQs4BBb/7dnig1FcmNG+AwBMOIYv+IDpQ8k5UACmRclQuMxEYEkYlNpDOAQU6Jc04o1dUIEsHQFW3IXo2IU3eANMeINd8IU46DPe8FWmlVIIVAAMEABMAFMt3EL2q0gZ+NI5jL0GjNJaRYAFYNRFXVQMRIEe8MrEtcejBQA8eD8VwgVaZMElpNwOsAC/C4AXQAAJLFRDPVQYbYATIlzf0AR0BcwmRAA50IHQhTJdOAMZYALYLQMZKAEVEABAyD0quwdcwIBbrEVTJQC85I1osAY8QNGKhb5FIFMeLIVSGAYFEAaAYSFc+NVgZcSYzE1J7AEmWNYWmAA2WAQ2iNZpLU5r9YFT/8xWV8THzqsF/8CDDyjXRYC9+bVOCnhY3kAHAaiGSVgGLzgGtzvPBthQVwWES9hJqAiAfO2NQIuDGf3T2wU7V1WCO1jfL5UAhf2CxZOAhFVYgx28NI2/t/wCC5jVHshY34hMJXVGL9XbCr6D8msyf7wEZcjGlFWGSPi0f6HehATRBnQBjajZfxXSSGjKJ+jZIy6AXHADR+QNGfU7TFCB56sEaKi+WrXiHH1BGHSDApDaLk6EJ4gFFbCAatjfcjiG/UXjSSgHL9hfZVBjLyiHSdhfTKgGTJDHciiHro2FXOAC2oyCuR0Bu93Cp1zRioSBAqhOHr6+WuUEIZCymx00FP/gPBawRxiwR2Xw0y94XN1gBSyg3E9+QQsYQQDQ3FeYS+b9QQ9YQ92jskBb1NJtQg4ITC4ggtWNPPiMAthlgl1+AjgVAGsQ1RXqjQi4AQSYzum0RSyoQN6AA9CsUehjABdY5C6YS1HwAEdWVAwoxEN81ut9RN3c3gK4gEpoATboxGgFxfI1xfMdReVUgReAgYuUgR64hOAIADwggPiFPUOEPRz4AGm4WVoAgDV+gNPzgsbUhRlKU39UOxpc0gDgR0FbgwamQWf0V6MyTAoeTQu2zyJwg4tEuoT14P8U4BNhvli1xhfwBqECGGsoAqZcBpHU27xdX4y1VIARaD/Fu0b/+LTWe4e66OHpm74fFoR3LKp78AYL0IIl6NHwOwQ3CFLeENonTkoJKAAqTgArzuqsnoMXPIQvZgFlKIdliOM0rgY4Rus1XmM0ZuM3juO1Tmu0Pmu1jus1xjw+4AMO9NQWLQAZ4NuYdYEq9gBNQOEpY91I5rwSKAOKLIERwIRdEMFNbgBWIIQlbMJP5tMvwIS7kwBOMOVC3cHT7AJqqEAoY13daOUGgGUuSMRIZYBaZtR/YYVc3uVd5gMmGIEvoIV/4Y160AQPMNf5RWZBsFkUcukiUIEDVAEi4Ocq1moEwEsibADe5QRJ9UQOENdG5I1fQIFjDQS/HucWMIXwRecN/1DnA2iHa3XnF5CBi3QDCahnpngDAlgEQ4y9+5ZfDIgGl60FACjolC1oEjw7NG1ib9A6rttJczyhBnbXrfPXRW0AaZjgD9joFq7hXCiAM3zFC/6CSyDpe4CDbPgPtkPRF8Bdo/oGl2ZKR5Bpv25vQ76DSxC93/AFWcVGIAgAMPyXU7iBwM4+7APRwV5GNF2DWlBqFniCRGhqIviAE/CXVGC+uWU/qy7JrbbiOdAGP1CBt45rtp5rNobjM37jMm7rs/5yMidzuv5ytT4Gui6HB8jjJFfyn52A2bPzwJ4+D8iEKTTsBV4DGkjsMphdDjRbhfWGOm0Af/gAy35CyiUCC/+wO83uAW14hVcg1NCmZhx4yE3rc2EeNEGA1NNlQtiW7sl+3QuoxFRngS9AhH8JtGigABBlSHMdgBtY3RNUBfp85g6APdlb5AQQgS64gTUc0m/AAE4I30UwBVMw50bsjdxEWBnYg3GuBAZg9vGFhi5Y5wNg5+QcgHd+8Q+I8f94AyJAdmS389hDAAxQ0Hso8mpQBpUNcLNb6CbuRbxDcF3gc4qOcrizVGk4Axj4ABkY+L6WgeQGgkPIzPGDgVd8AQ8PQ1kERxr8gmPAgzQodRTyBiBgcZHMgfYuvr6mcBhAgQFGoUsQyZTHcR3vDR73cesDcqK+aX+5hCiOww5wSe//OwQiWOJ/4cWKRkoVYOqSzFFtOIQdeHNlmMe0bvO6luswZ/Ood3o3n/q6bnq79gKlH+s1ngIWSAQu2ADAHlNO2ILYLksVCjRAt+TFpl0WKII30M8AILxhpgBGn9QJIAKK/QIQyGBosHTQ1sEuSAAcmPvRHULfAHXXDszXXt1Sn20ZeIJUR3W3l/Gi+oEbyGrrCwV1v4EIQNNpqAX6TG4wRdfY4wQ8pz4RoADdnTJtBk7wbfYT4A1oBwF4roQCqIRK6ETx3QAXmNZXqNYDUO8bAAEQMD6/HncDBgEisHMPVUiiYPcFhoNLiOkVT1kSTAVL5Q1duIQi2GwRZLsA2E7f/2DwKB/wo46GgP+ALXbx98ZGXp/O7nPRO0CBNfwpWaSF/3BoOLhZgLjXYI03IAa1aMnhxk2BhgxlfEABpwHFimsuAdECRIXGABPXUPyBA1WoUApOlkTlQUjFlg3s4OG4pECHmjULEPmgA+SaVAEuCbj0JUeOJTLYQGMTC8iDcl6cQj1Wblk5qU+vlptUFRMATOWqgn1K9emxali9KLuqbOzatFOhjn2LVmzaapMAAOjBJamLvh48cMIw0aW9gRVp9JBRQkYZJmVYFHnz5Ys3OxUjEOAygMEEzpwLFCnyBcSXWNAcdBHloJQD1F0S3IhGsV7FR4YLU9yymQsHBgx4E/+Q0gA3RVZRmFxAjvxJDzyI4NCmKCzU6wQoXSCgwIqiQDuXLBQBEl7CBASLzi/qG8pFKAzTDIN8tIUBBzac2JjCL+cERVooXlgQhQyVXFBJJbPYx8YGLmywwSs+HKDBARNCWAoOLwTCEEN34BHJJQGAIIcLnPRVYnqLYMDTPWvgYZAjQLz4AAABoLPGN4ZRBAkeL0wGwBcCACCAKi7FEUkARwogQBwUgVQRN3XIUICGUhbQg0EdMLDIAAMQQUQBH7wASUX1pAEIINk0YmSS3sAhEHcDFYSQFlPkAAMLdwSihA4v0KADIrg0QBtuFymjUQ5aqCCAZbg1g4NJJ0GqgEr/LOFYEUwSFHWBTTUl0kEBOjSwIjoBCEBqTDmMUAIlKrg1F1RnvWoWJlY59cBT1bwalVm5YhWXWLwCCytWk9iFFwBu3OfCIh6gOFhLxFH0S2JlKMYYC1/sIgAe1lhGEWZcdBYuZx+MVgQIRbihQGuqseYabO+FGp1t8QW6xhZcMIBAb74xQMAJaxB3jx3HJVfwEyyA4EsaTa6xQgKoOZCAdaEsskVFAqXyhQQbbyxDvuilV6ILYUxUmG33bIEAA5wswsYinHCwXz1r+AeggAYa2ILOH4ShhM84iBLhhAdAKAoCL7zQ0AcF3EGDhwG84EdfqLBXtbIpDjRNGru4aBAQ/8vgEUA2awgEEsa0IGKNKtegw801ccjG5BpFHokkIBRB+2SUSzPU0B0WANEByFvKQYQniIxZZiPFRNJ4AJGM3VLZcSJUVEOHFIA5AUufkQp8TGJkKKKKDkdRBR48ap11knoAqksg6YIHpktouulNoK6YDalJYpIDC0+oUU5TDyhDfFNUIb9WNcrEYkFYuQKQbZBvALCrsK+uletd1Zc1CSaTKFOWVHHh6mux2wNgDCecMEtB3NG5FG0PjlVbRglASPZFLd02IEVm4oaLXCAY4BfcMAfViKIUClRNxCgwGNtQZF4NgGA0MMAFBKjMN/giwr/cFCpdnEE5FxjhBRCmsP/amCE1qzFBdRBAqVA1IBUo4JgEZpKlEplCZC4EickmKAh8LSI/QhyAcBoQgf9Y4AUwwNkeZlGflpHIQRKSEIUOIApOSCBpXyoADFDgjbC9YAChgEYoSFIS9lSsSfWQxhsy4kaDfIFGbYKhQHQggTtszCChwQM3LtaANBjJSEeKA0huVJE0nKFvl2sIDFQQOJGdZ0sf4A9FtJamxjXOG5GoEZMM840AHCQhM6EJKT1VgM75sT9FEF0OBMATiiDBA5BSnQKs44EiQtAwqQABpkpQO9sdQglko1mSBPAGFcRiCsKbgvGKp4xyOJN4U5hCCRIRvLgkD5qwyqZTitfN5DX/BS3H86ZUcFUNrnCFenjJVql8EYBivDMSxYiDLtIQhzTQggCcQAABtlOpJl1mftQqgWPuR5pdVKYiC5ADuPgVLjeMZoBFKMAcWjOOUmigFAxMwAoGQxwJ0mZmC4tGGqQBB5OmAQ7RmMaNmoSLKDyhYBfYQwktsAtCUsQZInBAAhNYii50AQdFhCEkXsACjsGgAKYImciUhQDXGTJQShhAZ+pTHzZwwXWIQOILSoCzSrRgFhtQUIM2YAIJteMAaZ2iB6KQNMwdwg0vCAAeBPACR5EEFQowCRot5qQ2ik4LyoijKgBKETgo4Q4wuMMdXiCB0ABAGmP6oyBLFYAlVaoB/9xAWg9e0Fm3ngFpWjgEe0jSl/PIgSUCmUYcHvc4TT6OkK8ECRwCEJ7KjbIDnSKl4TxHkajSAhOhTNRHpCPLk9DSlrj04y5ZYDk/dAC6A6gJEc7AE1okCQCxGMEOyqFMZjLTm8abZiwMYYAZCE+83hRnN8O53mi+5Xhwae9Uolm8BwwPv+JNr/HSC02qlMVYhEDADU4xm8/hrQGQEJAMmODgMjRSMrvgVkWQIAcEdMY3nRmAJ/AwQPAcwgSq0YAoMnrRiK2gNio+cD1wQYAM7osLnCAA4qLaAFyEUKbJYYEFUIDZBiShCxjVgA9EMQ6gFpiODTiBUSUAAyd3gH0iW/9PX4TaySYJQQ6bWRkHYJZV2mz1BSow6hPs1AM3TGCsZXWBCSCU1jdHKBRu5a1ctSWAM3ChjHuFFEkqdjFrWCAhgmYVYRlGETtA6QMweHIWX4AH/tEGkKWyLGZfeY9UCKghi/QSC7SQiA1ISlJUHoAgxtTaurk2ErL9nB0CgAllZMQKOShApzjVASJ04A6+hSFFVAEAGBmklWmwiCZkKbHkKqB1EazIjViBhzdgwgJugC61qVsHkEwDu4FgQSCUAd4HgNfb4IbmA1TABwPkYgTktm8z213fdrNbvcOTN3+Lp0z4jhfc42ZmepdRLB+54QYRAAn8AFqYojKGCQ1mQiP/LfCGCd9IIBZuKL8YwGEPg8ACXyCAiDFa4hKzhqMV+ehkG3AKAvCLAyr3DQfjh2MRjvAJJehxHylCAVGUWAMkzmgX3HOxNZzAySx4sgw6sCCqrSfpLhjAv0rHEyEQQcsDQMAFMViHaKwhzGNmAYEM1IEWaENBLoCGWdGq1rNrQAGNxQlNwPSTAEQBAZGCVEk44Vc4qYAoWpCArIHwI1o0yU2s8ATfCiADRuNBspVsQGsnPcgrUyQOgUjqBzDnqQ64wbmVAPVJ9NpnrDUgGtYoJqpVbdgb2SESADjGAxyRkAJUwna41rVFKqIK4b4ICMK2yBZEUMvfr04BCEDcBJnd/wBaqIAFS/BlC/ww3eZDNwwLgwMtApHMKXjbu/r+9neZZ4hgqIHfxFv3ut1NvGrsoivkjze8+wvuERiCD4HYfvZHYH/vZv/bwnNKsSwQHIIHSvEBVCq8QMI5mIOpgMOhwDXkkiZsWYxZ3BnggQVknAUQQcfpXAYmkMi9ybIdmMmhnMqZwsrNmJi4BI7F1EyREAz0GGadAjXs3BSRWAKUWgA2AGLBwOEdXgEMgHq4ANJVzQ2Y4LLZgw5gwR18AAZQwAcQAAHcgBDcyFZFQRJx3Ve1ABuQFdmd1dlNSFr5QAI01iF0gBgeQhTYmScsAnIB30l4wN19Qy28AFHIYQ4AQf9dAZ4H3QMkEALbaRoM9MAlwEsDvEfjJQmpNEIhtUQcKNHSNMTluQGmFMAGINt6EMBgREMABEmQTJrpQd43NAKQHMMyZIQMiKHtYN4QtsTtAVtGCMCw8cQWIFcCmEACVEcCIAAlBUwD0IAEKB8LFMAE+MEEdMAA+AF0EcIpzAwKbBcQTNMUzMk0gZu4fdcUGIIhqNu96Zu9kVt4jV+9fcUUjEArUIIyaZ+97cAI5AB4fWMwoIEhUEEw7MB3ReMIBAMViAMVjAD37dvwOEVXEMJOTJYEvQcrFGBjHCATJCAILCBACcID0odvyIESXMKHWYAcvALOZaDO4VwCYEAqFd//4tXDKdzAynDZItAHARiYBzUAK5xBTKXgCM0cCKQCSFSACOic0GSgCAwVRehCHSxNlERJl3yAJyiBIOiAUeqAFEgBNxRGYTSJFDRiB0wAVU3ABCjBe6jCf2xdJeyBgVBCC3BAWWmhLIhCAohAKJylCPyFG0QBGd5aD0QPANwBJ8wB8EkMG7phLWDKHNLhjxTWilzG0lxeQxweHjgLSBBiMQECQDWJIiJh39jEI86aJK6hpNyA4rECCqgAJvyI4y1mBw4EIGQX+ABBUm0KtX0A8bkEJKwSMyIEAOiCJ2FALZkAC7GQLNqiCUKLLjrZ8j0BLyQCL0QBCtDACSDCCcwk/xyQQw9YQDNOATNO05xIo7flQLp9l3dhpzyqIwvMgBqMWyDQYzVagiHgH3iBYzVOQXdNwQx0AhpUARqggSXwQviNgHXWpzsCgyTcgiRUwQjsmzSO21dUQ/qMgWEJoCC+BAqUAEEtHBPkAAWiADrMi704JL9EZC2gAAoMkDhc5JBpYFl2JGjm0nuE5EiqHBtwwAhyAgWkJI6cwjM8QQG85AWwIAhw0gp0wU1qQDvo3DB4ACoqWOURAGEKDirolUkcaUncgG85JUWcgGBGl1ROpQ68BySgQCCoQBT0AOx5ZSUwQBaaFYQMDU4mwAdEgc8U5RlIIB4cCyeozhwcWy25wP8WNIkd1MIbPNtobAT+CEAxkI1FnAAB4Bqusd0HXAJAvYcuYGIxCcAhVgprgUAP5GBDJAJNSGYkHhtuWgcCRIC3IM0X4MElfEhsrcF7vFI0AAKSAMkDSMATJEKtoSYlucQuHcqhaAEA1FwDfMMKiEACvMIrdAEL/WpuJpjZ8CYMGMVXssAIqAGzqgA4joAxBEIPjMCzPqtzOmO2MiMzskArQON1MtMOxKN3wV8w5GMwGEJ7VgEVDEEVVEH4NSO6GgIamCs7wud7UgEaDME2AIO8fh985mt+SkIfhEAfSAIwGEM0OiezXqfw5IIgGGhhCIRAwAEKsMDQycATMMHBvID/QuJUbmRQxcWMDkxkBXIBC3WBA8jCMGiULDRQk5Dc4pncSLIMfqAoB3zAdqzWQJyCJ6Rg19HomNXINNxAzuEkieFA3HCHDuCaTfzikc4dXwkG5C0ZIUDm1zWfDtBGVgKIZ32VgSBIg0ADm4np0ECIBiQAIUQBEUDXTUTGFyANUurA3NLtCZyAHQiELlhsUfiO7+xAttQCdNgg03aAHGzKlyBCVCHm7kxaIzhLSMUBL00qrVlqD0xmps6icjmpJ5iZIx3DjxwibTAmHMRBHABCI5CKBZRAVFJbAchqS6SCBeSArCEEJuzaNFCAxATr7gJrAuCACebSiqBAD5SAUYAV/xesirNOgQqoQfPSpxo8a/jBq3NCJzjywfSWww6ogLsGwxQYgzuiQb7iKzAUAjJcwRCQwTOA57zma/uG7/tSAbtKQhM0wRDErzuua/hWwRAUwhUogiL8wR/sJzDkY3rCn3xawgyEWzmoAQsogzJUDwCIayAEQgw0SRrgwQgs32I02BJ0rI9VRCooYRNuDgEQAgWEgXECSBJxgizEYEaWZQiM3Ioh6MzqS32YAsxwAiFYxs6uQc+SEIHQVCO9QGFJgRngADUkMQ7gwA3cAAVsAbyYjRAQozC2gFSiQl0GH6S4AOi9UtX2TaVSFwq8RyrswgCJWYF06QSYwoJAAzS02f+YDg3asuUw2jFoSAYB1NKx1WIChILF5C0IKN8SLEEv7gD1BC5AfQPUSWWUGm5qqmQDiKax4EUkDFvBpcEMTWqUWGoN0cSWDMAN5MQHYAEGUGnVGp4bLIEEiAcAeMMaiC4MkW4kpMnuFIEERIlu1cQAEIDr6CoMpcIxFQHgAAEAoAOz5S4tAtUyv8YN+FMuDYTF2s+AcIEfcMEsMMMhGIMVOCv0Ni8f8MEUhF/0Um8zqoB1TtMINAE5NIEkUAH4uusQSIJ+3gLBNoEi8Cf8uqd7VsE8yzM998EttHP8xm/4SsIQKMIVXAEY1HMfOHQfjEET0GsnvPMQpED75qMjTFP/IMyA/QUDHwSDMVTBGOhC4L3EJeSd8pVBY7DAB8eBm7iYynCASfZGzNAAHCbRC3DCMGQkFGhgAlhMSKkYtuXIDfDGl1rVDluGBK2kJwRxgQTtC9RCNGRCjt7k2aKtJtTeI2CAZ1SlH5gCnGZqpLShRawBT5yA1TZEJdBEIhwCDZRxyVqACjyBgXQlWInVBmhh2XbhhCSAJ1hAIwtjATgcJhDBHMzi7t6mH2cCMAtyIUM2C+CPc8BBSw2EIBiuME7XdH0AJHhQYaRC9dzFXVhyAGJbJjsZDLgBJx+CDEAim8mibb6GCNBp/3yAp8TVk/GIn8ZyYcABIFjDJZHKrykW/+seAkBWSlEtAd/mQBHQQm0k8+4yM2woHjTDwRmwAGMMSFVWJWdUMxeIgx9YZ/PmQneKc/OKM7ZOUzBUwS0I9C2EQBOwAyMwQiEAsACHgHsT7EMXrEMXbD33934HuEDjMxn8gX7md8EqeEA79ALogi6MQRUAw/7Kg/0S9Dun9wjMgCHwQsA2wRhUtmk7XQA4Y1EsaBlIAIS+NEWkwkjSB8yY5Iz9Qi1knGPt9DiMg45GiAaIgFZ3EuTByw8YtW+g6CJ0WRjYBrQMHlQDLQvgwU3DAQXoHI+qFZU7gZh4kD9QACc8JGegggnAQ23e5eoggFYLRJMCnVrDHuUWAB6AhP9P4MFoWAAfFMhdh1VSvHECDIMcr1XaRoFUBqMfFAD+fIE4ILZtOoBsh4KPx5AFKF/xFi9kuFPgCoRtPEIdZHYLCKMwfsCQzLCv2cUx3IVH2KAgxoEm52CUuEEuuHYOyIAp1KZiz7ZfScEhXLEpHZ4F1MKfAhTpFoNwkwomqICTcfKtCdOPN4AqdNUSlEEh6/pZN8A7uILuCusywwbWOR1FRMMZLMZK/+IENBQXcAFw2h84Lm8stKshQGv8FTAQTO8IPMMYjIGC/0E+JAMU0MEqHMEq5EEyKHQh5AEUMIIt2IANmEHBdkMIdEMfuEM3jMEoLMACgAMP8MAmJLw9MwL/FEBBHnB8HpAAIwQ8I9iALdhCOCRDPCiCwbozQQeBuZ6jO6ZABmRAOuCA56zIbJXOJ2XE7BJyCagAnvrCis+skVsV0dMYjSeRBLgAT+/oFO24ArAEbeSSZQf5kNOHynUZFtBLRSw50BIIC0r1KeCAD5hdO/DoOFBAbHqQFNyAy7DMCD5MopeCmJO5HsCQBN1DWvcNW2NOAdDA4k7PDvgSTRlIIqRZWek5F6KdnwN6VR4CBRaBH9CiCSS6a7DQolfEL6jAgkJ6CbDAIYcqHJw1SJwCFlRxoBMjISheKgLAWnzPjFxyRUTDqae2DHAyF2GKxyQ25QOVxPjVAhDAdAmj/ylFwZB40FmnAepGAmxFApCMhwS4QYyekoHG0LJHugoAHkX4ww1Qe7C6CwHALI7oQhQwKHJU5Sx0xjUzAycMwRCIAy9YAjAAw772wTMYgxq4IxVQQvcyLEBMmTKCHDgeunhIi7AphBMcOPIgK3RlSJV4UFY0WLMGlx1WHhHqYiUS18gIJ3kc1GVnUzIoJPJMRLatULJwaxo0WOdkFA9wTYBREUoFzQg0QagAS2GJqSWhaKqIawIOJ057Db4FKOJIi5YcS5aosPBlVxycDX7cYLDIFBu2HBZ9UEUrEIgXPTYM06DhAF+/GkLpaFCvwaOchQ9PyxnhBhcGDDhAfhym6v/hBrg8Xaikec9mGCpeXFrgoe+Bdqb7dtGU095ZYTjYtGXDRlu6UqIc5HaQIIGCBDikHDZ8+AShArkKVCpwqEABPDh1RRIwHRMLJns0V6LUYkP3DQmGHRAv/rSGBISiFPDTYYKfQxZAFBmQoMsrB110m+hyRQjxKCUAXAJAFnZ4A49L4MgJp1MwGMCPCSAcYIIBCDHLsjVo+QKIB5RZRpkAErRsmjhQkAAGGGSQobkCPsuhhAlMoA+/LrrQDwOcFiCivfbW6+AORBpQjLB7GogjkgCOTDIAAb4owgIVWIChgA/OCFHBBlh5AYYSygBQBVoO+wEH3mqs8b4uEqDAMsv/UvlPhjKYKIALxyZggM4BlIADHWMIGWEKFabIRSpgggpqqBH8VGOKGZ6JASEeFog0hgVSAqmjR3TpSFOPcOmUlZJA/VRUhHA5yNRRwqHAhiGuMCOcELqhFKFUYrhFEiqQEgopYIJIQRIDxBliiFW2IWejwwhjTSNvlHEECEessCIHFQy8JA0iG2CMg23Z4IATyDBgRZUXnuwhFFH2Ku2vwAZbE9sgF7thlsdMkYwBTxK86jDMNMulkn/3+OwFPLboorTy9hIhAmUvywQDCii4YQAOTHlFg3Fuk+VM3m6A5DB9NYrAuEQKIJnkAmiA7sjpABihBCY006yF2Lqbo5Tx/8jr67z0OmDPPfjkM0E3B0rJjUYP+svphB66lKEEp1l4o9oQcWpmCwowIOADAigggAAMUrkSJ0QsyAGIDT9M8KwgASnxxBQLcINFFbRYwg8T9MMvN/1WwAkJOSaEcAL2CAGSsCGLVDKAxa1JIxo44Fgjcsij0cjynHB5wWkmuJTAl8OawSHGMvWDB00KzhouJ0juKOEJJmCekwMuZmdgQiHWyCYKN3pQYwQ1AB3hCBIkGYLQoZwKJpCBqiBnjDG6eV76MRZwVNROSbpe+1BDJfUjHjotSZcFpi+/jz4kITQIpJAyIIUMZlCjlTxEwU0UEYRZU/Wr1vDGgrO1YAWvAP8BAAKohZW0RbO2eIsQ0kgFuV7AglDshS8+UJcP2EWYtSkmJxyUAg4ew4B62YkLnljbvjLzLxUGTAVRQMENHOADvojHL2awQ06wxQO1cMIU3oGGXiiIrvtw7BQfs5w9EGGcDhRgiSdDAU7SIJ3pCEAFL5PBEzRTgBcAIg1w0IEIcIYa86BHSkz8GQgsgAATFI2NRDsaEojDAj5wqQx1HMEX3vAFBFlGEHLw4wDkAMgbyAEL0kjWYX6hgiXkQA1nE0CCONiAaLTNRChSkYpg8L8ldCABectPF1DXACEArk4QetAHgJSTZK0hDkta3CsX94VjAGAZ/5NAD14gjTU1wA7/mivDm2TgucNIwQmvyBvpuqCAGynrLIi4gwwuALsLzGIWtXvMBLighDUUIxCxiIXvgDeFYFiCVwYwwBBSYM4hUKF4kjBEMIwxhl84Iwb0jEFKSAU+8G1vn6XqHg/scJAI3DMk+gxoqSBFvunVKn1UMIBD33c8NPiOGcMAonkyoT/h5IQWdOuKABv5BQPCAVsfZAAPN2AKTngLC3DQBRpfcAcFyNAv6gIMHDUSyUieRQg4QAADEMCJn3IBAVjAxeUw54nkcMYzLXyBB/hympyBsgH3WIO+IHEDTrjABd1BhQI0UJ527MUBojhd5a50GEgoMRFLXOIhdKAYOxxpSQKw/8AS6ijNSsyCDV1VgCzCOJ4uECIQKkBRIkhmASepMTf2G5oHgqMRHbzsaXAqQ9TyuMfDaEIOXBiA7TyLADytCScRkAALcpADLQBBAGmAV07s0LYenOhEbsDkWIBQgDnISDc0ckXlNPHZUtpuAmA7zNoAUVcBuHJxADgGJpZRhCKA5gXc2OUjULA52LGABsP0gJlm5AD9KPOEh0FELGAmzTo9JjKgzVMtQGAMPoATUYYIQlAMEIT8GkAp5gQGMv4whkn9Qp+s6CcPDFyqBOvTnwVmsIMRfNAHN1h8I1lAEyQRLEkUIgX4DYIl+DACK/DCYujaSxe2oFGrcFQFagCpFv8aCYAAFGMN2NIBDjigQB5yog52SAUKLPACN8yBpurqCwaVgKx2XYUwV/mGELCGASxIGQNhwAISbmiYs/BLhSqUQQvvMIeojkcDPhDBaoiUrA9ulQ2ogAYqxIyPg7VjHLjpAgZ2ahkeKLFnh+hAJQ7xgsqloRGw3MFX8AonJrSghxuYgwPCeJp2DPYMRZCABOTmhi98AQSMJVpZb5MbyOYEDmeQARNOferLvgEEX/AFSQ+TiQEgoE5E/awfkrzLX8x2BKjNAR5cG0lWWCMSR/JG4+CQhi4GAAg50C1vjdaFGxhGEMK1k+0YYNy09k8ABZwikgIgS0wcQ7qKFXRaC4P/gi3BjgncPQwSQnGfoYk3mVsoL1ZogN5oYmdekWkvUOsgDfj2IBeI8t0MmLJf/eoXGAoPyhUkEQODsILiCLY4xSk8YQcrmMGfOnDGS5VPAxsYHBuWxH0dSoVg+C4XdDAxTbswiLOseMUNoEUPUistGD9AxjS2MY5jM5tuMaAOcGCFDl4g5AT4QIbjseBeQnGGsyhGMYbRYE40seNFxIYTcxIEzZOanS5/uQcEeIUFpVoaanisgzlBAgLY4NUNwNkHp0F7XzRQijvn+TB7ZmLPmJiIQA+60K/8ggq+woJEJ2IWpnABKiCNM0l3AQsvOMbZonSH6XxBjRoTxW1u0wVR/3jgBDmRRhRkwAd2c24EO2g1grC1hi1Y+5oMkINgdrk0p5VgCSz4gi4ulApvaEkGtP2ADD4AgxcoQwsy8A2NcqN3B+CgiLPHdu0JwYqqXm4NAZjELAso4yN9QRlAiG4RgFAEFLhWf+p2HRPm+ESs/7Wsnx4HjUKBgRAdbjA0cEN6L+AC6iQyFiGEGIAcWKEWLCAQKCHERmAGOsEAyInhymnh+EvhDGAiZMVURM7iOO4DPRB8dGETwmEUFmATFkDCFuwULg6gLM4dGGGdFo5XLKEo1IAPtGEYmI6C2qEUXOG4GgBkhkMVeoD3ciBacsARZAwQrionegoyOICrXECotP9JF5JOyEzg6VCjPHzABTyB/a5CMYgkkhogEziBE9iAEzZgNuxEm4LwcrgsOf4lF4KpB7ig6XLmYigArSwnGrIu7h5v7kwAHyRNjDTArLaA/yrDHiBBCqRAB05AB2gAEnUAEo4qihZnuZoEUKalBwzLD7YFFV7hACwIZ3zgzlAAAL6gli5tOvDA0z4v78ahrKih9BogDaIA/lZPBnqA1fToWhSEAhxDhB7DMQjAFtdkaditBGAABIDvuK4hErTEtgrgklhEsZoPFRIAHoTGjWSB+hpgCxzjp4qRAQihiNYEDvCAQ75vEgroSIpAGXag/KSrCIAN3daABgDkdVBN/sr/UAQ+LyAd4P6SaZmwAllQIBaeoACw6AkmYFsoZlseAwtU4RIWMBcc0L6KwhAabn0YDgMtcAa3wQncwVQMDCFGzsFSciVVUp+8ByVNxQ50wR2uoBAeCiSDoihErAXOrqb2QhRuYObeMK1UwRO4pPdSSwuWsMaccABoJ8fQkAMQAHekAele4AOysDTyUAO0wRPiQFkQhwy3AA1dIO7ibhEQINf4JyceIYXmsBLo0LBCQSvFCMUqgzC+YSzjbu4EcQvJbC8SYDWM6Cwi4AP8jAg6ADEPgQDOQJeMJBMFAA+azQqWgDJ77xAeYwNMgC4lTRQwIBWdC/0sAEnwYEwaqxQO/3EWx4EaFsYeUuEOmIAfYSeY0AgEfAEYL0MY2ascCcBjKmMx7uAJVE0GXuAZNQIOrCEAtEQ4q3FFMon5SuA7zMRoZMEDmqEBMIAcQ+insm/7DkMaQGC1HuAB3HG5tOJs0C89v4D91uYbaqEIUwTVQOAsMiEBYhFd6ic3QuHr0O0bEhJmArAAHnKluqVeOKFwLDIWcsEKRqAVKAFRZsCcJLThKPQCKzQk+SsokCEPwGAMUoIDTTJEYbKgRvRDEcIZ/uAKII5QQBIDbXAE+GAVwmPMKAgH0KrmEKMBVAE2maCOwMIKMCEAvvIbckIJJOQxCHQRuEAHJEcH7OIDLIYz8f+OE9yAxiyH6l4rJ/SSqzagq0wBAXDvhFiBHJ4AOeASLp9AAnIhAUhxPOxOBCLrSk7hA7iUL0URNSRPZ3Cq7QiTABCzA3qECIhACQivGOhKMqOlMsEiB9xgTjghC2dIjESBAmgAAJyLlr7AGwChFgZgDvCjFEoBYzBGFHBgYb4hApTgLu5CBXqgByTAAuCDBrghzU6BAAzQXowLZIBTNpngBcLmEdZgGuCAFpTTGlVEbjKpHOqGDeYAb6LPAapTCuCAAsjR3x6DEG7oXRqAG15AAlRrQ7xAxvBABYDAls4GCL7gK5HKPRGPS1CtSnJiBbpgGFATP3HDAUJBE+7NP1X/7wKwqACqiQFm4VsgkgBoYBcwkgUeEFFGYJzMKZ346wb+IByagAIqtglSRRzCIcM4FhhuJQWyQBGawBZC4A/IwAlsIAQ2kERBtKBSYgzIoCYdqiMvEEMr1CkMbgZ4IR5qCmE0wAPQESdUZzhSgRzcQDjnqAxyYAcCgAmrotqcspogcgCCww6s8hCiNO0QhkpTZvsIA0utTi+7FBq6Ay1x7yqsCks84QnOtDMqIU39ALAilYY84KiOKFsIoCzJ1s3mIB3w1E37Ak536TAigAAAtQNa4HCJ4AyA7zFfCQCAIFoS1QpaCHA4gMgitYLGgVIt1VKP4QsiIQ1U4Qa0sRs//29UEQAEDgQF/q8AALAEegBWQQAFroFIs0UtCHAtJlL7tLUBfgEEPDF4QUAVtu8eWkk55WYh5aY5MgkT6oYDOklo9AZfNeEUNCEMPsAwl4MQMEAQFmZNdAEF8EB1d6HbZAwAJEAFyFUCgIBcLeAaquJYvsEaiqBuBKQEAoH95HUYZGEYVoELtkEWcCNfhTIn/DMWTg1mciER7qAOHFgQ6kAQwkAQyOEQQmwGFnYGItR9zsm/CCACcOERTuER3oGEH6EZmkEPVFgP6IGF9WAFnEARQsAWRnaGa5hkZ1gRwAAMbOBVViAcdjgZ2MEGyAAHiviIjRgHxEEcaNacPlK/LP+hFQZCfrSh6e6uHcbKHNiOLTeqAVLBGBryAk5tCUaTCRVEE/zgQdZrW+Sg9NYABZIOa0sxjC5mAHqABoj0XRRDaAdDbLvKS5d0cFkhChYyZv4FBt4AAeY4Z4DyhIhECm7AO/hSASLvb9/0ey9kdQx3cBJ3PRY3FR5zuVjGKyS3MnPAAg7hIefgomzqBlAgDgAhlmM5DqYhFfJWARRAPwKyFIaBEwIBE3ZABbAoAIm5BF6gNkHAF/EgED6LAOHiMeqgcohkbU4gOAMQi3oATAjjEaxhOtLjZFaERUDAea2AAZpVeuVNAbz3BqqVNz1GW/PtaQCEkXjuC1yVffEZCF7/wBqwFCe+4RpoSX0v7QwshAJeYRjmgAsoYaFrozqTxjuxBAS06wIANscWqFvYgBkKrgRcZmE7gRfSKZ2GwL8koQl+4BH84QdW2IVbuKVZuAboIRNepQlm2IZJloZv+oZrGgzMIAlceKVXmh5cAQcaTkKNer+oIH4QhRdWAQ9Rw4LM7Hv5D4dy4osvADuiiXNUQADMWCMEIY0hhAvWq40bAA5OoFuJIIYsuS9EYRFy4QWsZJecDAPQ0Du4SqiQ0TJYYW0LgJj/pfhmaq3vjLRECQe6g2zJtllrxJhk4RW6QATgQQRGjbDRggAeJI0Rt2fOoBZcaYq6bTIXyZRzq05s/wY1KahNtaEHPPcLLBVEToFaXSAUeKOxyooTVEAZBuICWoGYKVr5ggxWC0RqWMAxTMFbnpkL7gAEBMA4ceIEYMBfo+kCSmA07QAOagEA3gAAWKBn2oqJmHecu2IWzlne8CMBMOAE1OIxFsFbTuoDish2c8L/YMZHWUApi4C2Lu3S9NkaxAYrGgEAHoArvuIFvnINMgEHPIAXLGGhKcESeGEOcAD31oQVQABAehRmHjI2tIE2mIEXNHgGSkCDjQKkzykFRNrEzykchKEZXLql6aGFayDGK+AHpuEUKkAKaIUhbECGc7rHbVgR2CEE7KACamAFasCn14Gl6YEayMBCj//avwzAEEQMRvcBc8MIqhMAp3DUdlkBCwoAOyghAPnA966hqtbg6JRACRwYC+oAC8JgC3zzrF8gre/OFDVgESoBrocyR9/wEegaEL2DDQYgr7EFM4YZO7AjFj4gHeq8TfHnDStjCxCgLA8bGkwgPOyOzJjOA2jgK6c5WDVZQkxpcPygB0R5OuoKco8wtKVFGWKhBcz5PtOlzDihB47h1sUNRFiBAgZgEWLbN/KmFGxbGSyABQIQ0SnamH/bAljtDXYgFiCjuIPuMWCgCMgCHSAnFbIhIY89AL8Mj6TmDcYCBg63Z5ZInCFXCyZgtzwpN9IEvSXDLQi2gSD6HvwPi2b/UwZyABNAoBqLL5gu7QVqYW38OQ4AwAvGEwi0AATU9QYUQKEXnMEpQVBCCamyRPHyatEGlgO0ocNngA8+PMRbgRcywMRTAJ1MHJ2GoHjIwBVcwQlg3gzMIAQ2IQZ+oAKSIIQfYedxoQKE4RT8ISWwAYhDoKZv2qaB3BZWYAUyIYRxYRM2IQJO4QRtwAlqshAkIetHmr8glhcMAIN9xxK0ARrSxRRJUTWuBGRs1w7IIQC3w9gpgQXwAH4XhBBI3WcgpDc14gSAN61riobYehES4QVca2iNyM/rWpJNAQcIPSf2upCxYzP4wA9Eoc7H6gA8YGFOyM8XYQPGfu4sfZHJ/6wvEAA+AkAVaoEGakFds0pwBCeN70CkTn2UFfUrKPMBeoA9UEEWTJuC9mIRouAYlmEZZEnGogESsmaQfMoDXACXE8CXAaDYA3AzAlTZAwFWxd3Z3eBbeIjrOGAWogYT3kD8gXkHRgBAN2MPvqwICgQEatMNLntwmsgNLGAZFL4Fdou38OMV5AAgXkxgQJANB04EsUhrcK/BGoc03FyYeIEJkyVFVHRIVECGGxYsJEi49NCewwb14giYtMzLA2Vf4jRocCOUuFyWKOncqdPSkF8PZ/6KUqJEmTIWW3BhNitRLD4zWkWdkStFBqtDrg4plOeKpAUxwsaIwCNCjB9lx/+WrSAM17tHcN/92ESWh127Y5zY4BF2VLcQgDeBtYt2U4V30U4JS8IXkt0YfMGFdWeD0apCkgzMGKGGTwtt0ERpENVlXJcuCVCL0DRzZkPXM3kQyDVixAwrfCjFwsPtJA9CE/wEHz7gQyqhIHoMUMA81BUPIuYkmKOAQYcouhqYnPmotclHGDix2UB+gws2OCK0Xo/L04VKF/a8v5CLCAIEOHB4oNYP+o1T2rWGzgt+jLcBNBuggooJPhzg4IMPDsPFDha8scMbILzxRgDFgOAHFwwMNEFwLcCAhwAopigAAEAs4eKLIyijQiIToCKLA6KINsxooiBgwTGYHFPNMQD/BJDGCQTIMcAABLngAnMmDPAGADuwMFEuFxQwUQkqWBCFBRbskOEOBXDCARumoMkBB1z0YMEXFe6ASZgjMDERfJUwoYIyF4L5ggVuiDhcBx08ocIDWmjRAjQKKoCKAtCEEsoAys1CkCkcLEKQG5ekoUsdGMSxBgpPZGnqBSVY8EIHfnRQQEcySHAHHg9191A9aaxUjRe8AiDTPTcksIo8vFCSU0475ZILH3IQcFwMRJUgw1FltMCLVHyUAFUwfFiSwT4ZhJsBP4y4s0AEYJ17rjNjtQsZWe+yhQtc2MCFi2HOLCBYuu408QcjITzGFw/d2GCGDTaEkwkPwghzyiO4/+CShDD+lDUwvBbb1c0VQxgzwwy8QCOLD1BocECDJmvQBQYPPfTNTHZsUQULS9Q2whKbUeLULtk9FAEFwwknXAeELNSAKiC8wIUGJrfzYMo9JnKHKgy11h13DYAnnnnkucDJDYis11p782EJXyJz+JDyAU5rMIwcF+7iSzEBvNEDF6AdmCA0rzQIoYNOyyIOhTsUHmbhO6jQAgMcEDQBAiPC8IWKKQIwxc0v1gwEmVyIjGMpopTCo4/LlF7EMUUEAEcEBCw5AAIMLOJCKKgkIAcAAhRh5Xx4sqCCCl+GmaEFuXCSJgeYmtlmmHHOucMIT+D5np7KMO8loBOYwgUXI/8SWsCeibYgXWomdFG+CQz0oFTjmGLKgBthGpPBLLzsAw0biVCSC55cqj9BC94rAAxggAI4BOhWuZpENSbRK5k8wgbC4scqkIGMFByLEsWiRCc0qCwuJCJbfGBCCyhRgo/NACqt6AS4spABFmYBAozY1wJmGAFnoCsGYDHLD8QSFrREoAKa8Ee9hvgIZwijLgMT2AJCsIIxxEAyd0EivE6BhCT44xFv+UEm1sEDH1qMLBWDRFhscIUqGCMWq9iRyQB3gNFQ4GqqoEAuemCz2mzmjq3gxQWegIKeNaAZBOBe0CbQAYXMRBV4UBrT2Pa0NoqiKXcI2xqCcjWrUYATnDj/zwbY4AJT3EA9WataA1jhHuntYQ8TeEUbT/YgH6QDfokjnArcwABTbJI8qODbGv9mslcQgHCGQ1ziJrCmNTluAm6YHIpwt0wgYO5FLAACJtwwCxc44HOhyyYOdlAEICyjCN800gluMAAcvG4Ai1iEBxYRikMIIABfYMETmCCf3r0AeGCSJSa6xM/fqSAQU6gQCAr3BjpFj3d6EhOFLBCIWXKhcQzYXnAOAQNlaMER4ksA+cx3mvR9yBSzWNMiODCLWNApBfuon0q3xw9ttKB/bhigBHrwgheAAAW1YIVD1gAHOEgDEADwwgIX6KsG4AKCeaAgMtqADAgggx+8AAZP/zbYCkq0oqr76MQMWFDCj6HBWy0M6zYycAQSNIGGC8jXDSOArhq2yyw6HMsCMnGKd+CCiLhAgjAsBhm7kAVjAvNrFC/GAykkwRlwwWIFMlGXCKSCL3BNyx84Bgw08IET81ilyYYxjG2IIxZ2tI1o72gbPuyDGYm4QCxQkIaTSEEOIQqRIAsZjZmkAg8W4MKOVukgk4kiD1yghBtOECCsNeQh76AAG8bDXK99ciYmeQ0pC1CJ/e2hEnvYgBpZ6SAfhKKhhAtTIHrAAvL2oAczvUMo/vYgpyXgA8IML4VGkD02LMJMbOJCMldEOSrdrAxLKEGA1QCAHhRgAF3AUY5Ah/8jKXWzCBAuggCiIQVyIuCci0BAOhdBiAAEAA8qMMo8KdKD3wUin2HqQYEOcqb7MqAFKrDQ4Qq6AwnwQXp5UgEQBgqmhrqBC/g9ph9iAQQrOCIRtdvo+ThxB+GEaE2Y4gIMEBeLlHJhCFyoH0pVSj9tgIYNXPBDqzrQgwAA4hpxSPM1rBHUlnhhEgAABBxSgYMEvGKCTW0DBPbM52ENgQoaxOA+rsoHqHzMELzIQFZamIVGF6LRoLjCGGaY1nS1VV1tNQtYkPCXMWSiGf646yNCPWrDePGvhIWMqvnKalTPtQK4CLVcaiAFZ4SAHd0IC1zDEg5GDGEIKaDCCKiwijn/cCEXM+iqCUsw2hkYwxApsEoWUEuJPfaxAS9bAGwdJ0g/1CEorBAACHS73QPMgxniCEU6/ECJJ9BAbN3pTkN+sAUKYIAChKCAvgmBgQh0Zxoo0c50q4vdSlRCAdtdWykGMIVgppgXy71lgmzkNPaaTAGxiKXDCxeIFthyuWciSAEmh7uSr6hKAU55CaYAAMWx4ZrZxNE1HQyEmkNYAGmoMDp3nuEMI8ATjWgEHoCQgyVYZI9PkMA9T8y8HcSiBWzgxCajbiY/HG7GdGqF9CjBhByEl6Eq+MAsDGIQks6iBYbKgRYoAQ2NcnTJTR4RMRkX0R5caAfVGMEQVrEKUPjd/+8TVLRKU5rBXOiPEoaoQhQCsYtdBAAAkygHr7xQpEhcAgcK0Gg6nNpUPvO5qchYBT/E0YlOpPCqhthHVhZ9FRdm4NGPzkMhBIOEGUqB0pduqw3PFYNe/yEcFbjiFev1lmYkQQqtHhhk0PIuVq/aLDFIBVl+MDEsRqwZK7AFO8JhFnbBdQFOQAawo22Jj3WCF5sZQQmZzS1L1C9ci+bHPhKxP2svpCFCGECQIxrmMwSFG5fwBgMwD+mwCrwAWlGxD+nwCn4AH0oAb61RD38kB1SXSZjEATggBTPxMg1hD6ngCdRlcAbXAunANGvDNAlwCJsDTDugYhGnN6gwB6XgN/+8dAChYHdN13Q70HHLtVxpQhCJYAEAMIQmxyI0I2ACxgIEZgEd8HLYJHMOMARv0E1AoALdJADSoAPk1HPopGH3cQaAEAcBsAyJon4WYShLx1D5FAsTEHWd1IOzcAhXR1BgogLRY3AXwHUqgAk8BnZu8AG54AZuEAuDGAsgoQJq9wRtlxoJAA+NaAKc4AbCMSIR5Th2VwTBlAtzkAegwImcSAeg0AudCHjDwgWWkAtX9TFqYAVqoAZT4IquOAWXowKllQu8UD/MsAraMEGitwrMwAzklxMZ1AnAkAVikAVj5Xrh4kKN1oyFQAKMMAqTtgC3d3v5olbqEgM2ZEOb4AT/TpAEP/AO/vAOxDcvzpBr7DJD3fAXfWALf6AIYEAKYGAERvAJn0AKpNAL94iPRjCP9kgKn0CP9BiQ//gJfXAW7QIW3XgFBhBtV5EChhAMI0AJ+wAuinaR4pIFQ3AEUFUAlICHBcBarSEIOIAQjcMmDOAHD8hTvhALuXA5VmBHMxAMvJAO80AHDXgBZwAHDdEQEmgS07AGJyAH56FJy7UINwAJa4AOu4ACILALIGCHlfCRH5kIsyALGtAOJ+gD0GB3d0dlXCBxCAINcyAa7cVIGuADnBAF8nU4FKICfnAmaXI8HNABKkCEeDCEK6I7Khdgd4kJh8ABCRZzonBNXAAC/w/2AkDwAp2ihV3IAF7IAOWkBGn2eA/gCDlgBVzFJV3CdITzBEC2CFFHdbOQC/LVJ4kTPfWXY0BgPVGgAgUwdmfSYmxyCClXCdBgAoyIGqjhAh/QAS0wItwTURMQY5jwlSrAAhlAB6D4iaPoiaNIAtJJQVlQCMBmAEEQDBLJGa44ArJ4OWrAGXcUDKWnE7zgfu5nLJRgABnQBvwAAfzQBkdwBI0WVssYVs1YnVlwBHRABgtQe5Q2Q9ioe24FFjaQD/pIkAK5oAzaoEZACg7Kj5+QoPY4oQBpj/3IoKTwBzmEQzgEfiQAbFcxohA5k2hgkRlJVmRADm6gP5VAXbkQkv/Z0RCCAGQsxgmzwAlcIA7GwBk+qgaxsJ5RFQwKKArDwIAG1wOt1QC3BQJPCQh2AAdCQIGZNB5OYgrioApwsAa64At9+AT7sz+VkAhssFtrMw6iMAB78pWFEwtc8ILkQZa7xUa9pQEIEAhtKUuFUwRg0qcUcpzV8AZfMCUnQiVHqHJ3CQBuwAGv8ISk4QA+0ppFIAGtiYWOmWGQiamTmQZp8Hi8UnNFxwIUkjQotgO5YKOjaQo66gaI45ZgkgMHhSdPMAJf95o/1oNzCVKJUAJMUAa4+Qrk44ioAQ0FwCrDIXd2+QbHiQnKqgKx8KJcwJyg0JzT+px+J53TiQyN9mv/BjAEBvCt4PqtwGAA49qtKQBsjfZUq+B5ngd6TiWf8kmfzYif+LmfWSAPWcAIV2Au03h7aJV7mLYAY0AKjPCP7MAOYOAEimADIdANY+AMdoANd/UN9CKOj4ANthCQAxkC9fII3aCx9cixsSaO/hBqJVsBK5AEN5SOJ7AATcAIY7VoLBQuELktvMAM21AIC9BTJ+AGL1pdWHIBrLUGMSAEN7A9ysIHrcAEmxEMM2AIVJAC4dqQlmAIXBAPOaIBCZCTTwACxQAIvhBeNMYCBSIezLVcftAlhMNjdvgeYio+atNGWjkaXXAIcnK3iJMLOcpJBiKnu2QyKCMKcqACeco8/1HgBwxAdmbLCX7QA19wISDwBbuAB1+gO0URYEWRA0RyNyYgc4VZCgnmIyIBBJT6AnhwDTqgJJjqhReGAzrAqd5QOUDCJwBAuX0KAmCSCwxgJmhiEJwwABm3cXTyrAVQT7P6dQ1FCG86l52kKbtaEbjpABulUQkQCsXqBwMgHAMwIlaHCYF6nIkjA7lwXXtwqvFAB9DpnJ4onXuGDPKqaN3akPL7rVJbvw2ZAo02n55HAhDAv/zLZ3q2VEcgBvNZn66Xn/lZCMiQDOGwCUgAoGg1oOmSkDbgBDFQMSaLDUN0V7E2ah7csUkwjwKpCN3wDXYVatiwDk5Aj4rgBAuARf9C5A+nULL+QA81YBbhIALe2AROQAYhcAUhep8HbEHayQfKoiw70QqoWHqoaAh84MSGALWWEG3yIC4XGW3Rdr9B0AmrIAulIDrDoAAdgF2G4qp6ygJQx7zLxQy8UKrMI5U/i0oMcoKjMQd34L1vUA14ewiJm0kuYB4xuEh0rAEOQASEm4PhNQJ+IHXNdSaNS2MZ8gZ4MIUgUQJcFWA5UA4CQCDlMw4OUAo4kmCcYAEioQKUKgGnqwPbu7qYygUD8LqduiJwNgkP8ACYsCIA4KTWw8dmwruY4gfGQGNmPAIskC0woC0sQKvW8ye3Kpdo4rwlAL0b4AAJdhqMaL2EQij/QdMBQggAedysXBXOlhwLPXAIdDAPf0etnAgK7NsGBNxo53qu8Wu/9IvFy5gFbaBn/bvP/rvPEKBn+XwE7juvB/x6zXgE8vCMVyAEtQeg/qouEuyh3RgOPDCONOzBwtfBw4cLPzAGDduwm4ANFj1q5CgXCwBr2CCO4ijSIl2ywiACHLoABeONOkwGTgAFJFDQhZABVZyM+jlW23CvGbANCW2vRD2f8ykGSj3ACDyzNDsE3jIHN5IjORIKMlAUJSABiNx0ZGtfvXs8ifA7bWmH1/UelTAL6RC3JjgaHkC4gfq9hZMIu5smfBuDZqpZGmAah3DIefo7cWmUG3AQjRte/046qJaL1QEmAZgAAMpABJ1bmJAtyi8gUxJgyl9gDUpgTj0XmQhwA68rhrgMeaLtYR/mzY9rAXLdy7PJAbyAg2tLOFFgxPTxHrPamkkDAj6mfyyGJghxCCVgNtNczRyVAAogB9lMBK0iZnI4hFOirCMg2/ARtCxwT7mwDekQD69QraDIznnQzvPZQvJsv94qtd4KbL+Wv0fAVHvWz+zdrvGqnzrtjMiYBVeQB7bwn/hNadcYsJkWAwbjDLEm0hqN0aOm0eTIwcKn0iOd0QlOw/7wAwtgBt2QLgsQDmbgjU5gBgcTDpWBDI/maE1trwiN0ARMwPMpnwQsn+6r4uk9wP8FjK9VnAUpsA0JQM2gDNmyYL1Ip9WFuwNN5tVziaNyKLzOOtvKol1MozajQcgDUDhvnceJg7icIJqiaQouMAdqZIJtNBoJAEtb/Za84MzHwwaDbQG3beZgwlXHjIQYsSJukBow98miHAh3cAczpSoogAiZ/Tqww7oDcAM0kAZiqJdEiDuR4A0BgCJ5WVBEUEuZchC7ewheqVCQmzguSR9gygfKrCq4PUv6FzuQTlKHwAJYQglOeE3DrQAf8AJF8AJwUgSR+wWE7s3VEAh8cCWzfQE0pQKHgKqhIAvYba3+y1QFLONGIM/mHc/lbRWvl96d197t/c//7L7HCOIFTZ//9PlodDB7lFYBtod7lZZ7zrAFTjAGNBzgwkfg6b7uGL3SFi3SJOvg/qDCEw6w+RIDK2DTTnAF3sgI8fDh9Imv2M6RLl7iAt3i7pzwYoAMYpDwSyXA7ssPR1AI/AAKnXtNqO4AjeoAnFAqTJB0cYIh8WUMi5y4s9nbBCVMYBILsz2mZck0cysaJkAAFqIh3uzNcAk7uyuXT7IjSr7WoiACd6CDNNYnFkAEObrba1LmDOWkpMpVV23JAgYEK3IHCnDxoAy6DuACUSCIdwAD5wUCNFAHS+JzXYgfN9Apg16E7wQIgBAJARAJywQCRAAiBEEQsFMAgVDzY4Ihb6AC4lsq/6Wi6aMaCKRKCEwSO4ofUaN+JxxAzYVJzaiRAAjQAYdABIewER2A+RIW2i0nA3tUAKWyR7teAHY/5aiPAKtwviTAzv8b0NYp48k++1YRzwet3vyc+/0s7QKc7fX54Qb9aNiODL1AAZNWe96u3+G+/BHQjSsgjjPs4Bosauxe/e4e7/LuD5ngBIIBsOhCabXXDYogAoyQDHohnfspD0ld8ASf4g2/VO/PVPKfz/n88PIv0BAgDm/wDKsAEKUcDHTQxcGrLq84yWDC5IkEC1/evAHxZofFHbH8cGLAiYNHBhMOXaS4o6IFC7EuULpQqUM6UeNEaYhZSoOCZ5h2SMQ08f9NlAFcGCDgWFQBTQ1Jx9EcVypUj4sWLFKkusMCkVkeF3Fgw4CDnB5fLIAIBOKFWQssSvApIaNEiRFABAB4scFEF4MDDYbyVIDIhw8wYLzAU2fAAASJES8mgCgNIAFz5wIAIKBYHMzZIgUIIACEHMRCGTDgwuWD1KgmqaqQ8cS1axkqvoAgW9vYgNG5R3M5xOJCSy54RTmIhzdBgkUdiBA51OHQcjd4IkemrALG6ycXXPd4YcHNhNEch5Im9CbQmxFD0oFahQwCsiNZCmXIkKL+kBT49edPYWRIliyOEKONNkiBgIQDE0QQQQjaaLANMeCLb75CAMygwgqPkEfDI/L/cGKMMRYQEQkRS1zghAUiSHHFGJxIhh12GIkxmXb0IcZGYohx5Qce/MHFH2z8eQdIIoMMMoZNuulmk3CcMENEFaNcwJkpTeyGHSds6QaJEG1g5AgwBRSTHzHbOAJCZAZEpo0113TwTQjifNNBUKrw6Q03QiloT4PwMoELGQLlI4c7LzL0DWP8GI0DBhbZ7YMdLqpI0pSya2mCdBwQxaZShhOFk0B6uhOAN+4obbzdEFBgU5k0sEmU4UKJYqJJqfIJBCJE48hRBnjpgaLazuqOhdZkYEsGFiyYywJO7sqroC4UIGS5AgoQ7AUa6sBhMQQW27axx6abDoAAskkDM8wA/9kMBQL8mGACBISagAs3pKLVJxTeSAu7C2JRAdizyrpDjsRIIw0BHHpzLRcuEBII2gS68GAAaonwqwBCpOtsOhVYiKW11/w9ixA/Ch4NgZDK82mXiQLpQRxt6LhiwgyyGCKDm2+2b2ecs7jwTPcUJGFBBeV8MMwJLawQwAwDzOKKPMJZIEQhTBRRihKlVDEcRshgRAQizDFHnXFsCEHEGGJYYJNRVgghnHBsCMeVFVYwI5l+oBgHS3b6eXIBtVWkUkWrR3GCnSa6WQAJLpHY5I88CgFTjDDNhPDyNglscHM4g44znVXkyCUQln0iJBS8UjeuiwQGKAEGtSTYgVQ87v+s6A5FheJCvAncuPXOSrXLhQNZNNW0U4PkAAETEFh2Hk8uwBMqMS5ULd5T4w/yACpbqaqIokOmN7h6IqCirayAQeih2CdKiIUFFSgrAoG76mc92mnlWA6wHlDwZNtubWtbhwEXZMQVmQAAIg0LRBcgvIGCDxDBD37gQmi4YIzvde8kHnPDE1ozGGCdDwSeIBhipNetQ/TANQUYQB76pLouuIBiFrPYIT5wBwFwJoeRSUssrtOaWIgMBImKVxHhNQBIrewNu4jC61gAPxVUQwCEUMAqVrGNQuTMZjijD30ydCYHFY1oRNvcmsRAuaQBiGlZ2IbTKpQHESguRCQikdX/BLeiCNggGeq4wdiSIYkmQMkZMRjkIAFnSEKqLZF4ZKSUqGS1FdjACU6wAYjW5jjHbcIVjPhEmSI0IFASSHNwctAVEAQKOsgsMZwozSHOcycqwnB1CvDDEp4IvzcAYBekKl1FiFg9lAllACq7E8tAEIvXJAIafBpHn/JwiDfMZiLOswDDTGiwAXBiDiZIwCuO083jKIATv7LV86iSi9AUkXyzEqGw1FesWKwFfpR5gQsU8E18KoAAcvDD/m74AiwA8DCgucEAbkABxwBiY+KKRBzgYIcFnisO10ABISJIBDmAZgB+uEPzlvhRavbADUG8DgxkgwIU0OYsniBCtyoY/70JDCAXIu2gHyIGw4iFYgDKKQABPlCAD0SBM0PlYQ+e+DE+yOAOYwHBMwjAHAIcIqoEyAUhpPI8JsLgfSyQQFim6AIPgDUUHvAAJ8qKAHHgYBvIwCIWj4AM97RhjEMTo9EINCAwOW2N8ghQXsGUDzBsYgxVo+PirlYirCHBCSIQmzpEoAhbbEKREVAkIil7yCg5Q2tVuiOKSlRY0Bp2E5gUrCbI0Au4vjVzbSpjnKy4nm0EIhBRkEP1SoODl37Aoz75gAJSd5eIhdMPt4TfLqazy13UbhfGIFj1wDOvYbJMIs5DwQ5Y0EE3dMC3fRIFXl6hgDuA9KNfCET4grKYCv8y4KZ44VMX8oCAWe3Co1ilyAe4hV4iREG+IDgDCtzZAxi4QQZu0Opg5gICBHzzfuGkQEaXc4hD3AGgAbzBDeRgYf19wDFx2FhnOhMJXcAhDQ+NaCqscYlL4AEPIJgNbShC3172wIc+dAMLSAcClPoXBVEgwAAHMEA/zDSIT0hEKIK74ASEAgHUsuEH3PCCAERiM5sJAAhUYNQ7sAAGd+gBbVCAhYyCxg8D0CgBrgrSKHjsDjAwqgVwMIc8oBIUeVgFnel8BX4goxBZxFBf4RqnBdF1aGQ02pqQlgW+VoivYdrQEQqBjDw0YRNrM2xhK3DYTYjgADcixjiS4YQQOMP/kJsldSNNfdjPVtqwY0CCEEjLNiGMohuMIAFc2YSMPCPDilfcRy5yEQsCu6EHEXlDDzR6mMUMs3keBYFFCUABAkQb2h+Idm+4WlwERia5u1hubZFdQTJjAQ/cFu8Igf2dUMzhngpOgAv0u2LncdsYEuTnsTdyZNXdZQ5cmJVyxVu6D2i0gi7N735xjOOzRCHAMpixhHUJAhys+zjwOE4olqM/IkSbEJ6gwA2i/WwMYAELGKjDFhKqQw8HoBEjhkPLXR4HGkThBXe4A2CWQ4AXvGHcAtj2uOUrUq3eIRbD3kWOU4qCM1SBzEsHjeiiQPNYHMLI+PRmAhSwZKgC5sne/5Ay1zdj5R5c2ag9iIKXebxRZDc9FxX5wrZ3EQiPabkHw/5CFRDmAQXk4Qp99lnf/yMf+TSaTYAe9KCLFqcHpRaNenVafCgnhg3R4UOjDe2lRXTpbsAjRzlSBzXGsekDsCMEf7CBGcKxgkmrTdSKBBwjB2e1VId2tKwe7SZizbZNOCGVyLATSCtiZRoX2A1ll0gUxDFmZJPZD7H4NwHuKYIEzOGbChCBxSXA1bC/wcPiWuIuo/n92oUfBD5PLm16cAc3uIET36Q466x+AxQkV+fbRkEV6u2HeutPVcdZsPsVAJb5Mq6eWyJCOLbky6/ZQIFAODocCwT0K7BYcDhuu/+Be3o+q6s+j5ODp9I4TyAAhOkWivG4aMMASHiMoaKyBNKFNYCDNZiGllsDXaiFF3iBM3g6NwAMQtgFX7iEbfOFnjMLTzg/GesyPMgxGkCpMyAEn1rCD6iCDyCEKAjCWCCCUKC+CrS6JMM6qQIMCZOyRoiEL4yEXbCAF1CBKIiCudOvIzyDfQozN9QtbhNAPHAZY5i7HjAGC9gFAnABs0IAD0gMHECYbdiGK8oiNboQ+VAtQBOaMUoQxLsrMxGDxptEpKEcSPuDBXC1qpmjErk0TwyHZBiHTksGV9gEKjlF1wMcJkmGF5kkudmESYM92COR2XOcwXIcIbC9UcA9J8j/A7j6RWQggVXAgWcAAQswBqFLxlg4D10yvvxzQ09oHvojACODPmu8QGgggK56gSj4F6LysOTqQDcMMyLwhHE7R7ezwQ/AO3xKAOjzAAzgNnQUAJQqQDfEv37aP+hrxyQjACLsOYDcBSzAqKYjMw2MgiI8QqPzLxkLuveJgrbbBTkIBRGwQnWgPg/wuIz7uI3zQBwYoAuLtg8gwXORMimLskgABBZkwTVYwTWQhlpAATyYwTN4AU+4A6HijB78QZtEQ58cPxo4wiPEgzOAtg0Uh48jAJe5STdAAIp8yuobKxy4OZ/6AE/QAS+0hjDEgyIYi+7oRhAIyl1QAkLIQALw/ziP+4D4GzcenMMoeIYeCMJnGAsC+EO7DMQfkwMsqAVVAARAiIO/9IVAqAJx2AZtWAUIWAV+eA8IMKXCE7Q4uYL3QJO3OrT4QBr4wLMsuoJ+2BJODC1ZhD0qkYJNoIBJMoO6qQFYUE1YWM3WdM3XbM0VgAVXmBtqSAYRYIQ6IwFaywPevALgBM48GE5GYATWOs73aI/XWoVQEIcqOA965DGMmk45EIf8kslphEorrD4R8ACc4w6wHCrxTDFx3CfqJACETC4a2DmWQUNj2EOK3E7qwwGE3MFt47mKMk8N1B8NdEru3E6K5IQUGr/ksk+25DYsOMt90k8CMEcaKDqhRP8BGlCfOuSyOkzPXRAHD+DOpxyrG6A2EH3CDkQYHCioCqMACiA5bjgXWmgEQHDRRmgEh2qANaDRloTBWlAxFUMpJVCCFzDJYggAXxAAXwiAbXsBsjvDKDgDAr2EoHxQskzKpCQEEFDS/9lQDxir7pRKaavKqwTDRqAFv2wEFYsmlaINFLsEHUjQDcy4jCOE+ONBOa1ST/BJY6DBuiSrQPzICiOAM2iEVEAXdIgDzRAX6cADzsADLKA2aRMHcbiBZ1CCQDiDQBgD2QoELDAGY/CEAnQCP9RTanAFV6AAuqGAFYAbEQiH2qM0EuHEWFyAdegGMzgcM3CFGlgB1WRN2Nz/1djs1UF4zUEIVjOggPjzBKSszo+kSDjKgwRg1jjTu0EsBCzCgUL4yCFAADIYAnHgAufU1BfATjbcQA3cSNI5UBqoy+5MV7LKUgT4ADOcwbHgDBSkMk9g1IwbV0I4AzwYUl/YVyPFgzPsQLLiTiwNBQLATiLlOfxUwmgb16f6ABzI0g4tWByAwkBQ2CHVQQHcMU/Ago7lVGPwWH190CcdSrIgu7nDSf3itrocK5clKwS4AUKggJm1KCyogx67gRJFSxQlBCWIA11Ig2sATKKNgxFrSRq10VTIhksIADxoS5SiARiVsloQUqstujOoQRpcwEvwBV+ggUs4ATVN0A+g/wAQpVksQDpu9ASdXVdqWNcS7VkCIISNowEvzIYxRbF+zRcco4EAuIRaoIEOBFEmhNNd6FojvQT/UlKXwVMPiNiP5FOPqwNr4AagTYNARQcUTLlIKIZaOIORm1nC7a+g/Fpf0AEMkJsVWIcKOIcKcIZzaAYpaIYKaIZzOAd6uNUVCNZB6Id+2MVNqBtJEgHfrdW6gYVfnc1f7dXYvNUaqAF6WIdz0AN6wFXZhAXlRV7tDVVy4DYegzajjNh1HV+ywoLD3cEiNa70RboabF9P+FYeZENGfTaNQwH0FdJdoIBPJd+3rVgafIGyAIEcmrIo44wkNFv61TglQFz05bm3i/8C5iLf8TVfIhVSBq4oajPKj8OCG5Dg8dXLskvcIr3fHazXj9PgfO3akjXdNQTg2iAdHawC8SVfHCAALCCEkRO5MOC4Cuth8KWAMFCCFZWov/xLaYCDaUjaG20AXXCgzvWGWvAGwKWFdHnRYrjiYvCFWvAFpNOx/kIBJw3cWjiBmKwDmsWAmkXjMPAvGmRDMohcOC7Rsp1ZkasDuwVDa/BLQKgFKmvapq2FYqAFWjgBJUBjQ6bjMKABElZc/vpfJmXDOD7Rg1ICa8CMoNUFwOxck0TJMKUFITiDMAgDkaNZQgiEJw1jXxCEG8gEYdADYagAT3SG2tWDGuBd3nWFQaD/hn7AZWroZVsO1t3dXe3N3tlcgSQQBtdthmb4AWdgZmZuhmZuZmWmhyRQXmEO1l3uL8Gk2RRF0Y98XHD2w48kBBog0q7t2n3t2l2g1Kxl50BI36KsWQTGYftl4PyFXHDG5xvwBB3DMRRASa/rOtBF4yfk5jDQAasl4XU+g2cgGHyGXDJQAi0eYQYGATQ2W4wGjDpo24d+3Bp+33+eaCHdYguuAyUsWwzAaCw4g3OmAURwaTKe0Jqc6axNZwzoaMglAFEOAwwI5TqoAww4KKFGUQzoaSGQBgbCjDSQhjg44iSuUXtoAKmOBsBsBK286kZYUVYg4hj13C1GASUA6y6m/wEx/oUxHmMlwIKd7mm1tmMdUNugLlG51lmP42lRFrkzkNoWzWO/LIbNgOIAqFoxNTFE0IFQVmvEDgM7FmktPsKwDuv+UgIKmGsfJgAMUIK/vNygjYNGKIYY/cIY/ctr0AEdyNqfDuWDPoGXFmOv1QHJZmVYju0kQN5bDlZXUId+oIYaSALd/eVgRV5hXoHotV3YhWbjdobjTm7kXm7ift3YFYZqDtUUVeQvy2E0rrC5jlydxQKynugtJumvhewuJt0tTuvQDbmQIwdF7tot9oW41lkcMAM+reE66OIcQ0la8MLNUII6UGy1Ru/6rgUB9+4d9K8wgO84xgEKUOTvZv/sNc1hHA45xUbwSMaBlf7WkQbcic7iS0jrQ37CnlaC745pRIhpte0vdtbBSzjwBC9RAhAEGA8DGFcCQdgCFL3xlC7qMEACiRpiOAgxFqyHpH0EqV4DiBLtBooDO1iDaBCxcxlTWoBiGtCBKUeBtyZrl0YEVfgFSDgBIdiC/q5xQZDxBX5rIUCBMOg4Nb8BVzgoCig5OA9iGigGb7DqRlCFMP3s/PYGaxBTy5WGE4DxOhCE0x50shbwLA5cK1/0xw7qs1RzHNeBOLDcSyZiPfZLo52ooCRtIehRGqdyVUAERDDrLV4AGnAHCqiBdRCGdaibQbhmV6AGWGjd2K4APaj/9QpYh9ylB1qnXdqVZVk27tlF7toldmB/3dp1btg9dlmugLoRhi0IhxPgYnIgh1DegjTvuB7u4TZP5C3G4l/w3Cw+XQVEgTMP68YeA9T26VAWBAafaBpIc26fdwoI67d+axTg40bIhs62amtw7UEvdDkX8AZPdJQ68G1nczYPg1oAXIKvhXCnASHw73UPgzNQgoRPeHGog7BGAXEHZF9IdLNWgopH7TrQgbI+65imgccWaxBAsVoQBG1P+HCggE6/eSXo9C1YAQzgeQzYgp/fAkGQdKNFapZjQSVugKhuyWiIqKBloKNtyZZjIECwhmsQdSqn8ietBS2HBFXw+gjQ/wEYFwQan3EheNIFQAFBSOkbx/EtuHlNuHkdoAXP5vdLf9EX5eumXmpEEIJO93Sy1wQaoHtaqIXCf+msn3IaGINbaHscp4AtkPShrXTMGFR0QZfNnqiJ4oZUuIbOh4RUUIVQ5/qYtHJ3cIUkSAJ6yAS7WYFXpnVcr3XWfX1bh2XXjf1j/3VkZ3ZklwJkh+Vmx/VMcIVWpodwEILApfFBl/GUHlUUdX5os2PDD+RAJvjCl9B7R4G0J+sT0AFyEITvF3SyRwTC53pfsPGDGtX0R9HIV3wJJesWjX9/d+2c93QaFwIyJnzqL/wjBAgMFAbeoFCwoBBaiGjRqtWwIQ0dYf/qhBFEzqIgIUoIGuxYkIISHTRoFCtJq9jJhohq6RBU8aVLQToc0vqlCpKqXwppjEGhw6fPWr5qbSTgsSMGVaq4pWLK7YSmLVKlasqkKaOUONLS6IIDZ83XNQ3EirU3tkE9sHCigVVLduyaaF7TxImDTtWJvDRO/LIJKRVgVakgSRGCRIgOIYqFLEB0Yi8NIVtWYMAwGQPlLYs3n2B4LRug0OiuAYpTunQcr3DspJKiA0nizTpVMdT5C/JjHb8kUu5deYtlHXGu1eVK13gc42mMK0WEKILjEzpOqIqTina2bOiasGNnwww1V5qSCBO2TliFdRXWr1e/Hr16+Onnu2f/b/++/XP499+vsSJTBehRsAUiNCihhCYIKgEcBQI52OCAJ6DEUDYP1bLSYxlCRkMt0ikhRIKCKCGiEg5VeCEiDD74oDsajnSCQ9bQAsiM11gjHWI5JqZbhT2qcmJElUH44BbULURLhSgVE5GITY6Y45AUrAAhZdONZGI2SqZES2JONilEZ7SogshNOdFGwwIR4XYhLQsINNCUA1kWQV5SnGDnAiBqsqcmICqGxAnH6ZLGV9OsMQ1aZ5kllqFkrfFoWHAxCmk0XF3TnCrQIQIYYLqkwgokEcA26mtSLKAQLXzpEFUmW7QqVSajIEHqAnllowoguKKTa3HJLWdHWHDo/xIBndKZaiqZd/WoUF4nOIaIFJr85yq1rQpywnDFDWqHcnAsRygr3qbRlCp34fWXNHAs4AQ7ivxhhhkrJDEvvfOet0587NWHHr968EsfwO3xp+9+9RmcRDhJ5LvCCs4uMOuOUUll2QrATSbIL5feujEt1tCmIV+P6YRIbIsltoAOCmWXKyKCWEzxy2DuldcvneEKWmjWAJJXrdPp4BoNM2ajsXYf6zDxZEljIEQEgynlI147moyYdBXDTHFwGSql1DW0KNsxjpspNt3WfwV2XXQgO6fK0b0p7WqooRIbgRRSIFHYrHaXGsG3XUUqVj0NCL7oWW+9JTjiiD8q13K6eP+aSgw3faoLK56ykkoEtdq5eV6Q4BQBJCcgocnoo/MpRN0naO7sXXcBgo51cQw6KKFsfeXV5aCfQDfdYppbrlI2kam76XzuuQnpJ3DDjbZcCbuaatOspdrslDueCTtg/PGHu4ooYkYmNSQhfjdJZGKvwv/Kly+/95r3Pr4Bzrc+wPnaL7/66yQxyAr34pvECgRBGNfYzVRVEYRVElgVMP1OWT9qznOeRR0xOWYBx7IgyiZoLoaMToEK3IIOyOQsm0SAFqmwzqXiAI6d0amFu3PWCZuSCnTQUCkRONp4kuCqTPBQCmf7kZjKRTcMEhBQv5ACDxPYqiVqIoJkSsU1Zrj/tUtlqoAoQ4wFIxBFTnHRhr+ATmfIhIhrQGUqS+ShJk4BCTWmgges+AHvpBDHCDQDdGnYShragijDFS5xfvxj4hy1OGFZBzDWoZw0WJFIwsytjhGAI6d4gLkC3q2SUqjA3OYmSXRIkZOHnJ1qIvWNuETjFKxQI+ia1slyASYGg3kl3WZVybzpQY6xS86gCqXHR63BDnE51KNG4R1bENMW23PXd/oBr27UoBvlE1+90kee8+DPffcij3nIkz5rtg9+3QwQN90njHCsIJvCUBgAqZEJYsmxnXiblWFmJQwkRAAcM6whJ+/ySlf+5S9LUUoMIPELz2HOc0qhYa7YNjoh/+gBCfOcpyZO4Dl+5sSQJ4RddTyXyriBTheyUyEKAUO3TSCBpKSbpxAgoUgozhCKNKRTO+/EO8KQrqalm+cCQnUTTkaRKT0VqUw5ZydVcqNyRn1c5CKQKYIKcXTC6BNUZ4ULXEgDF3bARTRwcYofnAJ0PwjVVk2ZBrbwUlKJ4iMg0wrIt4zyG3BgRRpYEQ254iKumDuFP3gQgbCq8pSs8McP5OgMujlDjs3gAVdB5w/A5DMV9rReVx7hlTWMUiz3eNQ06sotuLKCKY3lJCskKUlT/qCwhW2GFFCL2gjEgBvVmR2hDlU4XlZ2DeFwgi1CUEzdEvO28WJm+MYXXPHVIP8TK2BHPkjRi2Q4oXz32kQ4tXnOFVBjEDU4p/6yu01vWhOd19Qfw7BLr3V0wxX9oMYKTFnIUFmwbhWo2yXl6CmmxK6lnRJtaC93OY7CUW6u5FQh3Rvf90rBGZjkImB44CnrcHJc1oHEDwbDxr/AdXb11UWo3mtBJCyAwKcYVAyt89i5yW2jpxAdJe3W4bpxSjAhbgrsmhKq3WWSxoiU6yPmKo1P/UWS/QQMOGKg4vfejcDRkCyw5DLVqZ7iEbhw8lSvGhaxDK6Ph1PcWQT3CEBuWXCjRNQ34DJKYGF1lDlmMi54gFe/SlKuikwzax/5gznD8RSnwIU/8lu5GHaKFXb/eMQvfVnZBhCutpK1aio8pehEs6LRiESsnOFI52b8RdEe3RZlFUXbbrCjmJ4Ox3fkRa/zNZO44xOu+FbATFuwoxf56AUU8vFqRYSgG+c85yaiiTBqVLcGm+hGrvUnXvEGmzz0EMYKzJAwetGjXjZYbi96YYZ+uMIVK2gGXvH6g2ZImtuPlPOiRRxDymm10X7dcyq4ylU171XBiX435ui4bTrSWwoqxQUr8I3v+Z7w0tY5Jb5DC5hE9u2jqZAGhL1db2Idea5FjZ3j1F3QprU7AoNt58Ij4Og917fja4wAYvUK4VMwGg5YtUNm7bBn/bqx0YkOVYHbudoISKDmL/hC/3JCE4AXvOAMOgiJDoIe9BOwIpABEAAAkC4AAQQAEFT+Ixzi0IhGRKLqR2/6owQHCAFMAgBeFwAg/CgWaeDh5kU4RtIF4A1ApAEQVw9AAC4RADwAIABPb8A1viCBF9T8DhK4wwsuQeW3pCEAAJjEJLygAgmwQAIwcLzjX3ANQBb+GMu4/AMAEHY/CgIBCFjEIlywCA8sghMI+IA0BHf3BqQCAECQQAFkUAA3zN4NbvDE5sfidqa7XgtaGIALQoEK4Stg+KEIBSf8UIAOFOAQy38+EZp/B0T8sRYqsEIOtJADIAj+G5FgOvgbkYY+IuEGCMCBB9Kv/kW8ABPaB4IjHv/wgGUAYfE1l4AMOrABVMxBAQn4///NwQ2knloJzjSgAAssQQkooAIWwRd4Xd3lEeIIARFMQAdYoAUqnwQs3dLhwQ0kQBeYgAN0wQiOYBd4gCYUYJZJgRxMABe44AQwwAD4gQ4Ejuo1QDSgAAwswRJgX/yBXdYdzikIHRHiwU9AwlikgTcAwOLJgOxNQAKIYCmIQilowBQ6gANQQDQkDisQAAN8IQdwACdwAQMQwQkITiqgQBFYQA88wQXsQQuEoSlwwCJwABuwQSiYgA9owAFogB9aYRcQwM3d3wuAwHIAQiN4AxbIASMOgBw4ohwQgRwQAhIqztFB4NI1nVpF3dT/WV0kBEAkxIHiNALSHd4kCIA1ABIrlF0RnF3aBYD4XYM3gB/cxV0AeMPdpcIX8FwPSEAvAp7g/VHhHZ4XLIP9Qd7jwYDkARIcBMDlYd4x5B6Vdd7oVaPoLQICYMD4qaIAvB4MlAAMsADgKQEKBEIqKM7uGZ4jaJ8fmAIqDB88Fl8osIHyRV/0FUAB3GM+Tl+WCY43qEAObF/2CR4cfN/RLV0kjN9bZAIOnJ8HNCQO4MANEIAFFEEOWIHvLcP81d/9OV4HuIALKID/AWACCCA3BBIg5WAClgDjLQELAEHSJV0ASKDgKAEBDMAAZGAHtEABvAAHIh0OJMArvEIXkCAW/xalBwiBCtogC+ZkDE7ABMwgCqxeDi5gGSyBBGgBEAhAIwxe4kACBRAAEUgiWcoBBkSA4MDBEqoAECyB7A3AHIigA1AhXZZCFm6hDeKCF4JhGJIhAZzhGqQhCFiABDzBE8ChHHKAKSwCG5gCNJiABozDH0qmKDgAReqdzb1AapiGNSyiI34mTj4iBpwj4jSj13VdJuYe1AFC1XkiLIqi6pHiaSadaiLOKr5AEQBBK6IdKIZG1U1dI4QGaXDD063BNcwdHoCAERohCiDC6jVA4SFeMS5eMiLjC6gCMzqjRmpkNGLZGmzB54Ge6Ime6WHAFgJSKmACELweEOSACljAJf/QACL8wjaORSNcXe9ZgR8EXzyiggIcnwsoH/M5H/NFX4G6AfU1ylgEgApoH0ACAR6sxvf9ZCTAAVwIzhZ4gEgmgP+JpALgwBcoQ0D6niM4Av3lQOPVHAwUgCnwJ0mWJA4QYAGqJANe5Ut+gdLN5NNpAiPKgR/4ASQSQQ/8JAAMAAgSJRYe5QnqgApSmQ484gsyQAzOoA5QpQ7IQAlcZQ+qAQA0AhwETnGegFhGIplKYhgUXQOopeu9Hv75wRyA4FxOYRWOIAXc3SNQwBcyQBiOYRmiZWCqIWEaJmIqph2awh2igh7yoWT6oV0SAW7y3AsEnTWYRiISAk5eKqYOACX/Jk4zdh1qMl1tciprUt0nlipsCg4pIt0kHAPYqWLZqQBuFsEy4CgsHh0eXB0t4qLicIM3XIIA4MElXII3III1EOcfxYEAeIGyGiMyWid2Qp12zt8DTEIjiF0YeN54cgJ5ZqOF9qPgoAMmqEAJFMATxF4BfEDtOWds1qJ6at9HviPx+efwucAAQF8+FkAiNB++ugENiB2DAuT74YFYuF2pwqKFPh0GhAKHAmCH3gAeiOhFZl/8qUFH1hyLuiMqLOz/fSgPqGADPAICMmAJjCxMfp2ODg4rWEMtDKs3rGwtCACOciAeGKkJiKBROoAJLOlSCo4QAClUSmlU+sFU+lE0/+jAHYCjSwbkMQRAt97gGkjBWEbiAJRlHZwnHFiDALRizeVfxtZsKchpZXYBBtwdLlAAGeppGOopEfipKgBqYb5hJejpHJpCizomZC6qDyyqZRbipC4PN8ABN1BdAFhqpmIqBpyC4nTq4QEAb4Yq4qRBIhasqSbO1qkqqzouKxgt3+XmMhwDq0bCJeDBF+ABHvyqLXpD0+IdAGjt3/1dD9DAcyLrMRQjs1ZnMr5AJfpRM2Ied1ZrIGVo6IEkSKYfAmBB6iaOKqjnEswePjLvByDoKLJre2qB/sVr8f2nAtDr8xEovkLfB5yh4NyD4FgfQAYk963FJ8LdJzqdH1GAwv+SpAL03w0IACbkQA9mnxY4gjfeHwsUAAMswjtuKADiQO6q1QE23gIm8BR4XekybeJswSM+IpB2gB8IqdL9alCGYFGWIFJKQZMKzpMOAAI8pQzS4OqxAg2AAAiowINqASYEQBxcmT0ggdQSwdROrRwogdViLevCQAf4ZxRiIV2O4BaQLQUgAF9ygtoCZtuu4Qu44R7ELaE25qFCJh9qwB62gwY4gKOCAOD14gt4g9R5w+DmpBlH5aUSAmmmJdctLgc6ruBALii6ZkJS7tK5se/6ESugwP3V324KQCSI7uiWLiHfYupeA/0WwQvYHzCugfgmDrIuw7JSZ7MqYypCK+//TmseGyAGkJ7wgmTpIUAYPKfgZAMmTAHslWu5oqvt1UJpfuLShai7bsDxXa+8KsAGWOCA3mu+EugHMKlljS8LZ99AroEScuDRdWUgue+LbiwBZK39Yp/vceQOpqgM/C9IFt/CzgEBo+Qf0WgCK2DJNnDqhsEFnrEfTEBPZuKvIkAUiqBc4uwJenAB2mDPOiXQToDQnvALYKkMlEEZsAALKAMMr940CILUdsANS2KVosUa8HButmUB0PL/jWBlVmYCFHHilO3ZhiEHqC3bqiELu2ElVAIXeDQV260GDEMfHoBkDsPegkB1SoAYp+8HiDBOIwBOayriql4aZEMtIrOX/5JyHEhuLXopOt4x2nFlomy00XZkK47u3IHAzQ0yB6IuJAfAF3zB/ioj9dkg4kTyM6LoDsKAWUce9QljACjDAwAB/R2DN/jRI3Ry8KLCJ4vy8SKON7jf8pZr8+Ij9KoeLBveMWACAHxA8IWCSPbf9ULDBBAB8+Ej83VAJRRoASiB6j3yJZTvgwqAt0woB4pflsEBBfjfm0bhxlJAANTvEkQzRuYADMhAbG/tBASvYi+sAngA+IL1NyOgBCTwb6vAA8rk08EBFqSzU+qzBb5ALYauO7+CzXJwF+AAPXusDuTkCEspFzgik+rxGfwzEzghyQpADPsRLtTBZyr0IxIBAf+k9VjMYiuuJ+y5ABDXrBCXQgKkYOJEwxHz5SKA9FgIJmFeANzOAkobKh4makv7YWU6qgX43ePRtNTB3U3rtIXntBpD8h1/HUJ+BSAV9S2Coog3wnmOBbKqatJtMuLkIITXHKw64K/y3FaTbiZi9eMSdg+/wFf7URwAgCRfXg443hLYro5npzIsQ/wBwTGk4tPhQid7AEjaNSqEHl6nVS0ogxbAHj76dbqqHhzUwtVxtVYSQWJfr0jKqzpH9vNN9vNVKVjoAjj4wgvcQQ+wwAjYeSC8QSCowJ6zcCCAwAL4Ag2ggy6gww14KG4nQChgQABYJFb2IEY6nhvMNv7FIOj/EV+HekB1G3AtvIAFeDoL94AFDDfTPV00YME5R6WqJ4IKXPAXIEBcEmU8FyUONIPHgjBOZjcMykG/6nE/lwETlAGWlsBWljcXYkCmRjAB5O4aLGF8v14BhJ5I2rcDfK0I0DOV8XdHpy0HEMAvoCEKDKYKkHQlTMAUtygnIGre+qFLa0CDe/odmPXjBcA1UJ0AEEAMft4AyKBOayqaNsA9IOuqIh5qVuhaHWctJjxSh/VBfp2KC07RtniEtyLM/h3PiS4AlK6Nx/HcZa0iq4AyXgLlNbzisYC8xztaGzn9vbXdhe/HUoAHaGvw0TeUF2/qPt2Va0Ff46Pz4SMhuPJY/xRkJnJ19ukf9nqoh6KCLjcvm+drIhxCLARCIFgACGACJkzCMhC8dCYewVcDwR9eNVTDDrBhLOSCODAAJ4QCNMyBC3iCN7yB/dovD1qBW8aebDvhBIRnACt2bm96Wk0DDUSBBbAwqOum0tVCt97DqSc3VOako5YiAHwBAwhlzpKg5U83+AISoiDOdZPwlPL6CX93CYQ3E2SpCnTp6kXAEZsxpn4AJAxeMaxuEUjA7Ed78I3kBjtAKCCB7mIAAnx0GP43BxDBt7NeuA++G75hHM4hFSf4Hi64u3Oxp4ejWffA2qXvIUwpAyAxhuMC5RJjMSorIHt44qTFcTJdwhvsaP8Lbvo6ri4YLcpHuOHrHeBVNY1vPA5O6Bfk5pwDxAtEDQgWbHBNAIBjy5apWCIDBow7MFjAEGiwIJwARZY9eABkmbc1awq+o+DBRUpULla6QFCHJEaCtYoAkVCgQCWcO90MJKgxgIAAmIDk0NLBRahQClApcOoUFYICHQq4cZOoUqICT0aomOTFS7mvk46NXWZ2UrW0Y8uWVVsN7Newk8pNmRHL2BsLDpcssZLDigQZBWQULjwBwaJFKZ8q8IBEJsFpDUjC2cViSQkJJTKrUAYAj1A4MaMR8jMB9QDUExK9OAYAdhEGCUyY6GLCQRcHtnH8oBwZoxDVDCYQZzBAziX/maxeFGYig0l0FQAakYzZQIocBAO2TxiAHIO0gmusAShSs8jNRZxYJqBt+1UoKRjhUGDAgcEiDovuE4lAMBUUQNjriScKuKAFDjjhgA1TNmADGhM0GMcHDQ4YRwMNHCDiBQsiiqgHbwCJJAA8CECAgcRQTIw7QlgxqBEAvIBrGbCESuO68awJiscAfGwEjt/WiMNHARISoJHIpHlBog8l6EGFIsyD4QMJJHjhBTxC8ybIgtJoxEiFgLDpIpmsOcaRZRxxJAcYIPowIgl8os+bL2B7TYBIcsSFgpRCYQlQlwTJ8TqatLhpJ60OKYCQOeEgUSiijCpgg8YSaAwVBjqg/yqWAj2bBFRQ31rrLLVKneRUt9ZSy4u1WoWrrFbB8qIhFvgoYYS+cpDgiUUJOyy/xZJayjEhgJOMMhowK6GEMpYoQ4UvEgLgki4bKE211Vbj8Bg7v1CBE9ts043cLnCA5NjghiuOXTkQybEBVs64Nbp6o7Vmsus0wQEBFLn7To46ojFIFfPSS+8D7hZBIBQPLu0iARxOqMegaDD4jgE2GORiAjlOAFBAC5pjopJKJtiPQVNcYAMVCS18OUMH5JDAww9DHDGoE1NceGHiEMDixZhipJUhWoWKI1+DyONRKB8DAMTaIYs8MkmZdNFhIojelACIYyxw44M77sDyC2m5tP+ugS+LPOY8CYqwJrIzQVpzM63hLJO+AL44BpO+jwkgx1P6TIolVFaKSpBjiylCixxwooqqQz5oNCNIhypKiwK0eQqVOZwyhykGCkjkiR5anQSTUGMli63WW20LVbRgb/WssmqssRxawwJLmRlaYaKvXnEqzI3EFEuJsYaNTTfZZTN7Nocipg2gyzVwweA0bVErwDU7AVDBhfduyw1ic0+JDN4GlFjXuI7fxYg55+rlI1pvvsFoCwQ4WXE75AYl+AtAqIlNCrAwBLhAAcQSgQLOhZFvYIAD/WIDfxDABgIM5BsBAgEIVCCDJ1QCQQxK2QY4EaEJHQBmGuKQBezWg6f/kchEKuLPDPuFBV2MpxGY8MIDOsKQo6VvDUExklCaFofrSE2IAECSkpj0oa15ZQduIMAH3GClInwBD9UiSGUaEYBIGOkLRbDAF+AmE28cAwgfcYRg3GCYN92BBpGJxkaUAQRHAEEZAgicK/zUFFT8KRQISBxwLqGMQ+FEK5ErwAd8soY0TA0TjctcpZ6SgM45RRt+YMEU5CIrV62lLGIZ1etcB0pTnqVGrEqL7uCSu9zxTgKxGN1OcKI/xSxmJaFYiSaYRxlfLKtZmYkeAKRFvYLgImHaUw33MFG2b7lAXF0olzRvcL5e1mN97Gqfu5bzAj7Uq145AIFIxrOGFaBE/zH94o4clIARWgTQJjYhAn9cgEsFuCdi1hzPxRRjCgUxiAi/ANmAVPCEC+CkBbPQ2AYcxDKXoRCF7dDQzFj4IU94wxowJIIMF2GK/NRwYDGJBFx4yMOzBMCIMtHIEInoo5RuMQ6QOhIgIsOciNhNBhJQwTK+RoQPhG1sWdJiQezQCG98MSFe+wJNzYTGZdiRjTJo49aUo9IA4NGOeNSjQQTXR13+CXHHugQQGofIWWrlA5ewziOFKKnMscEplnwKJxJhAVfOiCx4JSUpT9XXT56FdqxTZe1idwxa5fWVu8tdNcrBgidoBSf5qedkCeeCQaZrDb98VrOaNcxiWisVFP/I3mqW+YJmNlMCEbrN+KRpm2r2sgHYHA4DtjmngsQPnEx4ggpAUAu0XcsVSkmJYrhDgPkY5J0CVIFNOoCi4zUlFCKImHiUhgEEcIAD/jSFKdhAhI/dI0ACAkEsLgDCDiiUQWxwgSlMOI4DtAOFGSqFHDrUxifI4A61yGiJNqoYD6wnnT8b2BaH0kOPPAAAKE2fRvCkRCMp2CAxFaKRmAq/F7gBBm3EMEQk8NQCDIAIknMDliyAhzQYBA6A2K8A8MA3PFAXIwF4qiO0YJPBSHUwEbkDCtB3VbL+WK0G+cENAOlHQAryWL4gq+Nmqci0kmQabDWSpKxQAE7MoSkKmAP/J3KhjK/gjpUzmksqEbtKUc6llagScyrDzGY2t1KxulOGXicxBRjkogAZm6ywNuACDwySYjKJyWUyw9kyuI2YCbaW4LKFGi6UtplhTC1upKmbV5TvBjBOl2y5wIBO09Z93fzmE+rVCgmAAHBcJTJTUBFgAnxsPIiAJ9eW0IEZCkspl7rBgPeZmJRNkBPeBRAN8LALEMCgvFOZwEId1J4MHcAHEdXAfF8Agg3jNwA74u8tObGI/6YzDLzWiDI68gBHeORvL0VxABo8RAh7yXJCqbBBdHHhDLtJqjDoMBA+TASfArUIJt5iA+AQh0aQSIhfCMCJA10Qbzz1qUW5MWGm/7pjIPp4TFpQRqoLAgki/3Epf2QJAniJvrHmgMmQKwARFkmDtU4tgJPiRAIVAI0OAOErD9gdmMlsWFQeFgB0UbOpSIXX2yHWCz5HumHFcledJzZ3ZFaGDLjQ58UIy88eCEP6hOTLHhS6DM1C9GcLkgoCZItjq/nAC8rWzB6EYly5IR9tboAL9P1mi5rAGKiJw00Lkxqcu0V1kAINCRxgyiUIoAC6Yl2EKC1XAh2g7fEKl0AKTGMyGbGufhqkH1MIew0a7JAMLlB6k2mMDWx40AZMUKED4AOFFaK2tXF8h0t4w0d4kMMtKVtPBIS7IHNUxkfUpKZJvBvFLcbEa2BjJP91pw3hPJp38F/wgQzL4AP53ncBOiYHlkvkBTqQBtpS3IguJnHhkQlAHcfEpsG4oSq/ssjFM/5jAVirARH4uFKYksBAllyl8KAoEKUDEoEqWK4A4qgBomzCvgUwLgCuoIELRmDOnk537irq1kzMygE2AADOXIkudifN2Gyx2izOMHB3LHCxJiHoVMAPHqT3PMADsAD/MCImfolZmqUMnGUHEq0WQOvsUKN9JmDtnAkE3u4V5E43xOUVMi22bBDvFlAQuODTaKvvEKHhCEJeAI8JLkC3eOsHG+AeCAIJQsE9oCIUug0D9IkyrEEAjgEOjyHyeAbrksIDMCDzeo3zuCv/uzyGMlRhg/aC9PagZFpAY1bGBTYAGhLAB6LtZVCoFAag2jQMvy5hR1hs93rPzxQDJn5D+NSE+B5gEgTg+X6ixfamA50vR9Ig+uQtMuzgwnCMEjssc/rH36wPS67hOqIhDgDh4BDuRtSvjmjsUN6vKrIvbHSgBinDx7TAGYHg/gyiGYJrKUAHDUkOONZAAFHucabCGz/A5SgjDmoB4bbRCphgFrQhF6Zgh3bOHTNQLJROVarhGOBRzcSCzMCM6e5Rd3QOd/hR5wIyBfFKLYIuFqpOZYbrDpcxCtegFnrA0Mogp6SE7AjiFIKQXdRujMqmCO5AAZKQXMjHBBKAAuzg/+6uox7qYDtoiwPYhQiw8O+6UCZ3Cw+ApCCmQRMUoDbOMBQUYw1RDAX2Ip5gwA+ChfI8oGEwQKUwgAuwS2NMoaP8cA0AUWQ6qLzKqwX8KfUaZAMSIEPawRElShQk0QKoiDBsD/cCAAV2TwZbYrgWYetuciOIL42UId2WkRuc6TXwhBQHrgHi4KiK5Gkio96yr40IoypgYBm04BCOA2B+amy4AcVU7BeLxBtOTCbWr8Zq7CHiD2xggBDuQAmqZzw24sdqbKgIohlwQJcaw/8QoJ0iwzIG8HE2ZSpCTAG/IQ72q0QsAOWeoAWeQBkykOfeMQTP7C1OULH40c12Byyibv8Z4FE5M1AFV4UFWdACBoA9AGwGGRIjEOHrdjDsDm0HWAwPfCvzzC4ji0M1PmAjvwAEPNIB5pM+W4skB4ZijigKp6EOqNAKaYsLXjIL4yUQSI3UvPAJaOYSMJMytsA9bsMEnMLPOrEgpAEEgADygAAGBuCWrs5PPGAL0mcLmjK7+HARpJIqX0AFyEsnKiFBGIATuKBfEEABnu0RNWAsaSb7zvL2fOQL5IA9kKclOBFt7EAA0iirOiLBSnEaruEStIRHelTdHCkSgBGlCLP6Ju79YICsCshfQMynPEEyK7QRfLFKncYmM9OQfkwNBEgArCENpCENRgNHfosZa6LGcgD/CKolD6Xg8IiFcwIpNsfDFBvHcQzQAA+BKhIQpmDOUPmABeZMOi2Q6ZwzBGukUg0rdfoKr+TxHS+wHaUTzMCiRp5OLsSiVYJOiV5AHIDN2wghaY5FFSBSBnawBHLKAswzDAkCEjDyOBBgArjADa4IBDChI+cgCR2gFJR1Pkfy8n6j4ew0JYHVCouDAdxlQJnDQEmvCxWUQethBbogCXfSkjjhfyo0KK3kStyAQ3lvMVACAUJUJrZgAO6DE7aLQfxwGlQhKFWU9ECoEnKhEp4ABOq0PioELC8EHyqEC2gm/ioR9wQABbRTJQJFMcIgSEhCGo70I9QIGp9mGddgNEZj/yRGllDSIDCdZvoIghuqDwY8Eye4lDH3ZxFUowPCtIwI4kvMr0rPNE1jbE2d8SHcQGw8wWiN9gUYtDTrDzXxrwL+1DWXAgF0AAoJDgVosxI2pQA74BAIgMca4BsAIUwE4FtGQAZY4AFc6QEqULGiU7FUgAXKAQOFzsF4JOgykEbWzG3LwW1r5FVE0B39MVQBVyxARVUtwA84ods8gBDwMwq/EyLFcweXwAKI6Qt8qyAigAC0iT0nwA3KBgTC6A7mgFlLwXTnE2IwgPCecOCu4xHCwD//M0Bh0iBYoUB1SyYvgGYEgEEfwRXoEzdG0jF0IEdaVgXU9SYmoEN7DzZHAv8jwqBeGWC7UE8OjosqVcAqK4EQEypYuUN/avRGoW0cECAKLCD+wqZHJVY7+yyXhosTOpEk0oBjkxQIEgxqohAOECFLsMhOQmNBlYYVrXRl46X64M+AE7MmrKyjvpQA7kAVDGJnD+4XI6EUCUIzyUoLOhMnPmAnZCAKlJbAxqT+gqwgkOBPL4VzFGBqgQMOOIgbEfVmI+drw5alvkANuKIc0jZtw2KHda4C/XYE4vZUk27orjPoTOVTizOxRFGJmvhInLgDjfg6VSnoWFCJLABIEwMDXoR5ZvVWb1UiKRcT3gAAMJcgIkAOuIM9iWMC7gB0wwgGSHdZ57hZE0B1n1D/PyuGELajX34VAeQgHGv3BbbVC3XXAv7XInFAFBxgkXcjQhHguAqCGzhIAg7lJtq19xYDB5aHdRtAEMSBtu5VK8WBaqeyXz3kKiuBF5ySu1RmDnxgHCQqoiqEfM2Xg6kID4oEBLgAUAwHkOopLlkWADaTxu7IfkNKSGggqNDjivAgDjAigJ2GgploRzc4Zs+jAPasZkGMkdDmSyJBgns2DqJmiy4h4oT2CVRuUT/AE0CYMiIBT38MD3LEhPvvnhoDB6hWSVz4JgxwU4jgZg8BBfIFTIboDWBgBg5s+HKY3PiWbXN4Ci6AD+RCUuMsb1EQo8Nib5XzLTrQwR5Mmosh/wCKIRKKoRFImqSzYYJ3gUM94AO4OF0ggVbLgAm+WAXG+Dyv4wTSmFoz8g5CFwT0wg3kuBREoahR146DZAwF7QkfARJO4ASkgAak4AR0oKpPIQ9JQl4KOXcV9JnP2AMWeY5tIwE8gPFiQhVU1EqW4CYYQBP9zAUGADJkQhCiF7sWhA0GQJ/Tei9YKJUrIb04YQM2oHNc70Y1AAF6wJYXyQ1yOShQAAc84HBE7k/e9zqkAQ8288fqF2S77h6U2UrG5DyOwZn98lEEODJa1ioWiSe4VAUoJSVURp1e7ToMrmcnuIKD6JwzeDAKYFHWWUzjpgjuSJ5zRBgOr5LuWYX1Wf8m0gAEcmAJHOeftdbfUMA6xFaIjGEEcjiNcti7d1hu6yIH1IASZqAa3FYFP9UC0zuj2/sEy0FS4dsLli91MMGjQToSACEO9jsKtJMC9GlAC8KLZaAEmEAideoLdiCnCyI71HgI3Rg+jdUNTCAJi/qocyOpC2KpMYJi/EEIBEEJQFzElUAIVAFecGGQc7dbD/mGCKICwtrClxViGgha0xp5JYAIpLcOJ0uvfyMPlQCU7wNl8nqvTxnZQEhgpZcNBNsFoGEOTgi+3CtDEtt8ecKxBQAEDsiXjQyYr4Mbhvk0x0TesvpaUEDf1PU8rggzYyKafSS/sXRH4e+WC0AFJsn/Yo/jBiI5bSa4Zyk4j9fAnMfEKB6CKhJp5QoguGUih2isuA1CGDzgKebgUlAYkoGDFXzTSqZCa/+ZCKybMsTWSFZ0B6ZgbUt9+BZ6h3dgBIwhF3JBbnsod9hbo11pb8FbscDb1lHwwMrtu+NbbRd6GZYPTwJgFw6BE/67lwacpiWyBKLlDRacILIDMTh3AjzhDeBTjCackUsBR8VamjAAJe9OcPxTRouDCwAZXrZaxQ35Esa0ATZBBIaB27k9N0xgAMYUrXtAXdmaCDgAef49JXocWShGCOQANe6aQQbAWKaSoFTgyC9AYGeBuwR7A0LhlS0EvuArQzhBsWmpsXWZ/5dDARr4T+TM9Tqu4Qs0u8bqVwAAAV7goInOHAheIOBA+FGc5mhS2xuMJDTyJA7SwBowwXFUwnBSYjuYuwFGpEqPSpwvDo2I8SF+2xtZLtExIugfQLPn2SA0AdLvedKdIp+BAxB8k601fdP9TQkmAw7cUADegAVUQIdJvbsPzLvLYQSCwRJyYQToftan8wTReyAFMtZrXW1LyiN4fYcOTPE9AgQLEjYCgQsIgPEa0iBSYaYNHHicHQ9o4ToavH2IYwCiAA++YIyK4ANsw3SnzahFAWLkddMaQHA8jSUBVA4g4cTP4EC7sPRo5sUKYgvindvlywESYNeUBhGiQAJYQP8C2NrWAP7f85xQCWIBgvA/a7ad6oFfqxLfWID7l21l+mwDXtm9ND6+OL7KWc4NQOASWOwFEGDkQ87/XMCyBfxbMGfllcjlMcIOlADDAAKGBAlAJBTBA6eBQoVwIgV4KCBAnIUK6zVI9aKHhDs97kTx5OmOihyVNqA6GcqFCwQ4hFCM8zCSzAAy46yhqHBNgGNAHGnRkkNGhwIdEg0dioUbToWAMD3oqQUIQoqaPChQkACrVgUIdOC82SANCAsWVBQg0qGDH7Vpz9yMZk0AgFgjpjywq+zug7zl9u4tF8uSgUB2+/L10rcc4geKGy9uzDhy3wfLEktmXPly3geROU//9muY814v1SYBOI3pEIEIS5emulNGRhkmJWir+AICD601FhvoGDCBQXAuwgdEwfPFAggQH0yU0vA8uigHXba0bn2KAgPiDDgw2E4E0VJcZ54weXIh/QUWFvDoWkihi6jnGqCXMkEBbE5EniSwkCBQB6aopBIqLhjoghxSLKTfAkT44ccEwX03gRI3qfKCBS+oAMMFBVxQSSUTmLIBGxtsAM0cPrRzgAYHsFhfKHdYQEQBNhYAwiUCXPICAtCEgooCQaKSkgd16JdNETkA8dOSQABwCSD63YTLCx/AIAMMAhk0FUVpQPSQRK2lAoIMMhTwxI0FuJFDDgVAMySQoXiA/4CFC8EUpkOReGPTUjodo8wyTQpFVKFD3aHUUtdgsgxUUiW0UCZWXRWKCFiFwpVLY4KgQqdPsJXWWh241cA0calgzA554aXXZqBNQYklwUwRGl+gLcNXZYjpWg6vl/WaWGaQKebZXbSKZpldxVoG7CRemCbAHQSccB1FqURRggy11bbEbSAAkM0a9yj02wDfCVfcC8hZ8EURBZjgwHzQQTddddXilB0DCCzCgXfgQTJeeUyol54E7b2nkCsO1KfBOBqIIkoCGOjXwDc03AEggDAMMKALKRkIshys5bSQFDoooYQggoRRxxaCILHGGqqgoCGHIIIoIokmoqjiOC+2eP+ADz5AI9IhZ9kIAkQ9QnOVkE2jYqR+tCgJRA5ARQWAAI1QfFEdBZhp5kAqdLnQl2FGNNFS3LzgxpkFJFKA0W6MVMBJT8+JgCDTNBAzIAFElGckfZLMdyQAHLOMT0F1UEkHaD1OSKI4NeUIEA9ERXYDSGBAAAWdd07BBx/UAfC4hKsy0hJLELVW62pFkZAdjYBwRyDl0GqX5azmftcIuRgygmZ+5WUrsIwhVg2jmJTDLLKRbbbMA154dvsIfBxrWDnKMK/98KBxhphpAARCCLX3NsANtrLRRlsOX7yBhyp8KyQEcAzMcn+6eOygnAWHODcvh5WiXtY5n0IgoR0G8Mv/XwggAMAY1ABWlEcGBLuABMbGCoVEwwyiYFh9BpiAAi5kGjpwg5aWoKURbeBAHmuhCxzYGlxcAxKqQAQkbnjDU+wNQzXr0B72EKIW6OxEKRLaz1gktFAQgkZHw5HSEBCkps1hSB4QBEVqUbWqXe1JWuMaDzyxpq9lCQYHgVTZwPSQtOGETGZS01Dm5iaTTLFpLvAAFhISM1oIICKAo0kappSTSMglcT4h1FEOgRTJUWRRT/HJoyiyhUllJQGUvEpXroM6CSxBAqxjix/Q4on3SCMSUejBFE6pF8tZzlaFGUEnRqCGznyPeLOM3gOqEQAAMI8xt3PeskTDmVWNIBid/+DDLlfVOyrMgHeWEQ1pJgFNCxBiAQaUxguyVRsm0EYCuMEDOihSvwnlbwIDUBf/knOIV8gigA8bRxfyIML5XSdf3enXuQigSIVUyTwVNNguEHYKD3RQAz5wWAcVoAmc4EIHWZKBBMw0AQKZg4UEguFShPCBQzzIDwMw1wCs2ABVjCVDHaoEECvRAg6U6EQb6NnPNNAOmCrADUwcyiFUsEcBRIETTFPAHJompCpeUUlXsxpOu4iTCBijAB+4kZYkkLmwgCkigGgNN0BgQhsN5UZ0C9JPsyIkFxACLGvQY9b4SJPByXMNjZCLFxzxACsYMi1oOUTkWrOoyl3ukQvZQv8oKElJEwA2ATgwHwQbUIse5EB1jXNd6zyRQTvUwhh1AcIUtGCXzD5FL9qbwgxeuQPv0XK0s+QlX8phveAli5fK4uwUgsEHQ7zSL3jZwQwMYQDgMUYZvLOcZyZxjEnswBjUpAjXGiAN9c1GBtvs5jcXUj/unGsCclAXbsaSiFdEh2EDLIW9DNgABH5nEQwwhb8IcI2AXWBgF9hDwSzwT4VEoB8dHIcP6uMwBegBJ49QwtfaZqYajU5ldWhZHTCwhR+0poQ1UouEGDAAO/FwQyU9aUo3wAkizgFoLGpHTA+QgA/UNBFEOCoAdjqkrwZpTgltQD3WgEWr5cAKS1JB1rb/Js8GRAALRgujmdRFsTV8aY9/C0BVlxIHFGjJjWsaiQw24NOmJSAUoaBABhsAh52ctcgSuUmQ/QaASURPCyVgXFrO3IEPpFdtRaicMoDwpDRQBAN/TYBgBQvYwh5WIYnV5Oo60IIODEAtDyIEwOqBgljsYAqWvYsjNMu7zPIhGKoqbWia17xTziAWlJgBpqcwAli+KhjBQIMhLDGCvmhWBbGlwhByMatiEa+XiZkEJu4whtZ4mSHXZJ82S2CQ3MhvIZro6Lm+w4UBoAAPY0kOEV6xsOd0sIMOeEU8j7uQUxDgXBwg73fwuZRTKMEYd3CDGy6QJoN9YdhISMBA2yFA/w14YEEUYQUY3SDGAphi34vwAA5YgoMbDIACD8xxCbXaAQlxwQ8WqkcqUACCDLEARBaexQa0oeEuvEIBOOh4wG8ghw+oIBFGOUsP8CAXT7ggypO8CtRAyrdLKKlNNNaCjQUgpRxHgBA16rGZ7kADrsEkp1RtTZKXfKOiFGAkT4Byy8FKgWgwZBdF+ALR02hGBvltkIkrgdHQnJYPDBsn17AAkxyJBzkvhM6BTUAXBqvn1iR2CSUoQQt44QfV6J0AWFgQHAJhjFNattGQbtUDrDeDHVxatJvlrQp2mdlAwNYQQehBLy1Xjh1YT9G4GwEaTG1qSxjTs8sEtSEMAQxgNP8BGIZQ1u7+0phJVMMCQTfuUqwpgbprkwllYEERhD1CQdjv2BPwgw6QAwIUvODZCxvowx72XQNGYNsM4ES37QlufKEgChboAQtK8H0JqCsVCsmEfOpzX4ZRoxk4gQQWiNBUty3iJB4jkjlSUuVT7PngREl4hBh+Ew9XMyzwBCYVRBaXYTxzX0ETNDGlASGmAg2GFlCVcis3SXMAVlDTYjGDCBaQAyPRJkBgAVkTCTfRGw1wAjz3NjbSVEDHNUOWU0ZmdChwBzDwNVrVZEvwZFqRABhoDgogDvoXQcuGcpfgDd4QCY3wR36ydYNUEAiHZmKHVyDAJFUIAGrHNxSAFXb/xoV4hgMjsxRzpzrtxQIsQAiB4AtxgA5xkBBpEAg9wFu9dFmFh0ypxT2kZSvbMwIzEDydB1vBYAm8gD3MM1yxYAi2g1q39XmLmAKzMgWGwAcjEAinZwi5IAm3cAtVAAyxtFmF8SuyFwVCcFy7hmUgsARlUBvM5VBF0B7k52WCkGzTJRxygAK0cAl4EABfkE7yIW3PRx3X1hoWAQnU1y/m5R0EIA0kcxOn0APoVkHsgQfk1wAY0AXDUB8H4DD1gQMFJ18qeIOVwAZEMiRCgn8UIIQGdwcItxYT0AENJ4ASdzMhIiIYpmELeAAM6CIQSAAEUCME4AZvIBd3AGVX8XQK/+ACgkBWqlBkeAAAcLYDN5Z1KPgBh7RVQHdYcUB0RYdkNAgD5oaDcPRkGDhYPiUHDwQH1hAT1xAHcZAGf4RtgCBIuTQJyrA6/ec4aXEI4oFkZhcVP/EFWNgAWkhJr2ACb/d2hAWGU4IIGkF3LUAJsDQCmscCuZALz7ALuxAIsSB4p8Roc3gXhHd4ywQamXc7clg9wLMDmhcMhlBqVJACwJBqhfFahhgMI/AGw2QIoPd5KZACrTACpxcMkmcIVIAGwCAJTdAHt7B6daEXhYcXXqAMseAOFHOCDAICubct2uR7uSGNfAOL34EA57JwKHAJY7EcciALz2GN00ZA4NUAP/9AffzCBt3GAB+QjBB0ClGQHh/iXuvxAiggP9NAARDTMAwzDqJwA+eoEFKASGmhVVE0jnGCAbeZYyeQjmliFAnXAV5xERBXFgRogCEyAfSogPd4jz7QIj4QYhagktwQB4DgDV9wGnewckAFVgoQCmEAFnCAAp2iAhckATlgAQKAB5EQkVIwkWhRKAVwB5eAZBmJVDgRB3hQgx/gNm+kAjrYUj0IWD4Vd/zxAi9QdZhgdUhFimsQB43gEAIwCQ+gAmlSFFGokxJqAUBhhWoUlFv4Cm5XlJQ0AEnJIHNXd4nAC1qpBmqgAlypBlOwpFy5lZj1lZnFWw8wA9dDW6zFAn3/+FqkJph5iQZVMARVUAWB9wA7IHl6WWp6+aVoYABDEKZ56aVoQJhUYJi30Ad32gTiwJirUg4zkAux8Dx3EQvksIReFjPyBAelWRY90AN11wPKgQdHxjdbgAADgACXygUIkGykuRwgEAVuQAAYgAE3wAmLsAj7MgBygATfcD43MYzfYQqLMJveEXUVMT88cAa7STAsoALA2QCPcAPygl8PIwquIHUUgQREMGiMYxTQ6TRxckd7dgKe4AZp8jaJMAFEwJ3oAHEZ0gMFiDMoxQYmog1FxCL36CIuMgeEoAKHoBpnQVMC8AZ3QAT7SAE3cK/5egOa8AgKkQb92SZLsFgf/0ig3iB1FmEROmCTznkIMHAJL7hHW4ZjC2ER3MCRbWMjcANHTLChI5kACEBviFCDdwBnynBWE4sTafCeMClIFvAET6BRaEYAM7pINbokPomjQsmjXdCjCXAD3MggNMACdFcGRJoII6ACSHqkTMq0TtqkmIVZg5dZQDADTIA7cah5VVCXU2CIi7immpgFTYCJVbBoI9AKoFcFi0iYnyemQyAJVCAJwCCnc0uYVUAFRwAGeXsFeQsGwEAYvWQ9vGAJgccqKgBLbxAIu4ACKDAGKCAEv7CfvlAEnRIFKvB9vtcekoMLNXQJNIAIl1ALoGsNtOCdINADDJAOXaC6spCaDv/gAIKFAYRTLbA5XhxgXuT1AVm3jHWQHu7Vmyzwm6qwBhEwqjdADTjgAR4gApVCAf0KTnLAjmc2AVEEVCsWCtEqu9YZRivYAYfAneDgnRYAnieFUiulgOf6UuopYmjmB2QEAF/wAZzwb/MLcALXYmEBAgMrsAI7ggJgoDghBAvrOERwBzSrEHHgEDTxEDknoRTakW5jI3OjoRi4hZPECZoisk8lActQBMdgogwCBykKCI0AEZiQLVDYvTTQGoBgdjcLBF8gqTlKSTxLw5SUnLq2C0NbBkuQCH7ADFyglUl6pEN8pFbAB0s7h5aFWY/2aIdXAmoghzsQC4RQBYGAl2r/+6XAEKaSQAZXAJd/6bWLmLZsCwyFMARkQAZDQAVpO6dyaghuK7Z2eqeZ6LdToHl8QAW8YABoQGldeXhL0CvQlJaBQMhw4GVwgAeGe4qxAX4iiAdqxAoUgADBEZrEwQVyQAO18AUvsMlcIAvxMm3FWQoJAHM5RhEWQbv1NKsMQAgR2QCnkKvq0ZsXBAK00ADCIALzAjGq+3YTgxOCwAvFF70T8FMESb2hYA762RrW+QT4xr0FwJ1pcIvLxjbhKa47U0Qugq7pKQLr60k09b6HQJA8WEmhgJD+mr+qs78fmDUGC8BogWZoQQgG3AAYeRpy4b+unAYU+lBnkiaH8AQZ/3oBcnQVHpO8OABSiEAI5iYQcHYMAICyCwEHIzwTf4MJLGCDC0sEKowT9zChX/AFJAoAkUoROkvDPSsHyinRKKDDRdsCfsAFbIBqU2AFQyzEauCXp6QGmPWkXakMe4g7t2MMTUAOkiCmX3sLhikJkqAIZJC3Q3ALcTrGX1sFBrDUTRDHTWDUbUwFVFAIyKAITRACidkHY62YVWB6XZ0BBkCYjvhofdp5VhwItwC5FAEHu1A1OVACs9HIrbgQuEAIoekvyIbJiLDJRRAFDDAMzjesovAKG2jKEJTK/TKbi8AFrXyCN8EKXsNelZAewFvLa5AEuUxQHiQKXaAJQYYBmf8KHA8mkjxIKS5wJMucjm5TCYXCnXEQutQsAwYIRCmFzSrSYS91ACJACCAQKmrhBkUQznMgkndWzjAnFvqrOgJasBGpBASQ3Gf2AfQcB2EG3vm8FPs8EFmiJhJcABxAIC7Qb8iLAwUUAaLzNTDQKVWHY1OyBiOsohBxDACCwkRwAoB0EVHQJjkgAVpQBI1wgiZdlCh9ZTjxDShQdzuMUuQ0AbPADIPLpFqwpEu61026lVLbaCrQCrmg01WpmJKQC2zslod5py8uCW5rtzPe1QYADFZ9mHKcmLcQt2K6xkud430gtmPdB+7QBwswBkcdBGjAl3MKPE18SsUEicHwDFX/rAuHSlZ4kNcjQHd9HY0LwQoY8B394h3eIQeIoMkiKgGKTR8eBB0JANnYhsrbxgVl3i+X7cqwnB6e7bu8CgK1sAZbkAcN82H1MQwJQG/7udqTzAARYgp3RsFNYw4ekNrSegfN7EYfkNvIxylM4NnhOQvBbUT3CCPFLXJpwY5+8AQj+AVEMFhvh2fLC3Nrs1h+xr8j7Q0RKQgPcmbL2t1LAQhhFlwkCCmGSt4AciZuA5KoAFjQPWXw3VSH0DYDYd+jSNEJLBcv0M9wQ1e1t0bavs5A0AglvYUnzbOvgIytwZ8TXgKVECESonDMMARPSRhHmlpKupUhrgKxUAWZGAz9/x4CTeC2bnuJdmqnRE7WWP0HWI3VmEjWBv/iWi0J4kDwYv3wL/7iC8AD4JCJa5wCa023W6tpfGAJgCkOVfALELQ3MQcENFYCXc4euQEO2fYBY25Px4gIiEAz3afYjN0iD5MAmmJ7yqhjBEAcdm7ZWBBkrxwFH2KAHgK8KIAIaxAf1whT6ecBQIsLCUQcE8AFG+DslYSfHsCdRC8F+Gbbb6PpB8yQ73NNny6Ps4Bx53tEQLOe6yho4PwFBICBsN6zU3a/cfAC1M2rD7kLAYBHObHrcqCdrYMFQJvfAOAFwWUa/2tcEzoQWtJGTfZQG9CFPRsKBXQCRuNzLAAERRAJe//zZY3A+ivakByS0QOsAwKOEba+JOOuQa5Q7g3OswmQ7kthBxK+1+3+7goHHETQA7HACzntO9ezpCNgBVwptZg1AlVg5GT9B4wABfkABcmQD4zADnkrCTbwBwtvCyGA8DoeAt3QB+xv5EY+BokZAg4/1vNv/7dgC3a6ADHAAwDBY5SkKimGZABGBY1CKjOmOJrCJ1gnS4bEAfPVYI1GjhsbNKilzIqWJUtKlGBhAQQeXR8b8KDAgQEHDotmMiACqRYICxZ6LBpWSsNQUUM1iBKh4+NGjy4/1msQgQCDCQxucuCCxanLU2cuXKj09cIeCXjw0FrjSpQPDe18HBg3FAf/t62nCMyySpUBtC4JTPhVkEDBYA9SnDaVcqfAkwKNCxxyg6LBvTQBBHz5oqJELrCVPM/StoETtDk+2h04reGAahEfVPjpMKGDnwIWAHwhksCviS68eScIpcSlrhc5RixhgTwHiACXAkRzCidMhwGxrfshBGnrGkAAvHiZBEBAADjb4+CRIAEGjCcyGrsBkkOGi929+5oIteWj1A4dGsuQQQULvJmGI5e4aySSSAJYUIAigFCvsUQ6IAKFplxK5QWTSspBhUg8iuaGwBKw7zcTKJCmo+FekKEEGcqopIUJZhxggha44OWQEaaYQo0pLKpixylG4MOYHXicAgg1tJhC/wVjxgjBnT6aSAaKKqG4AoIrGCEhjzySicfKZKpMxolu+kDzzDOldGeTGHhYAE00/wAjHyigsPNOPcUc84pCJGniFkmoYKgTQ5AMxhBLUshgGzLQuUfFjQrU6BJltCApB5NGwOSLS1Jx6QcKrFqkVJoYIECVnXrqgZNhijJqNQ2GSWqprW49YaqZZpFJJiwu3OiUKAoAa4+w9mDhBRBqScUMWFdrZ6hSbkgjUo9OuYEDThiwiQNUHIDHARP+SmAOwgw70KUT3CiA3cY+aFepBioTAAAALGDhK88+22ADbUgzDTWB20rgAwtgk20CN2zDTbcS7QNOCJfA0TC5EkzKwf82PLwpz6VowiACYepmuwPUw7rz4phJVg4A2DXiuCS99QB8z4IcyjDFLxJNVEC/BnLtr78n3Ei2kVvXgAMQBZcOIABMIJQAwEMKqLBjA1mJQoLkluiwEY8eEdFh3/pKgALomBoOhJPKKCFGLmbkgotcYlFhx0CGHCGXIZowZscRYmkoEIiASLJHY3yJAcoxFrDhzjy2IWEVx7cZogoymljHmQqc2WQBzxeIAfQ3ebBDF10S7+PMPpywMx8SkKGDjlW2kZwRZ845Z506/7iliSEWWsiQYHYIhA8qgrBkBENSEAeFX8DhQZeNrF0qJC2AsMKKkiT44o1L6ProBwK2lan/W1StoQUFVl2FVYO4iFIA3Qu3+3kqLqzqlQGtbmXFK7Au4EwlWCCgTzlhKONYDVw00AUKpKsBzsABB0yhLQ6wYQ4O6ALEdCMYBKALV4phjGPaRYOP0Kte+NKXsfYwAVNsgA2kacsBZJiaA7RGBf2RTQsM9oUiEOEvvREXxEIhsY+oIgomYcHFSpCx25DHKdHAgh+qMwE/UNEPWDCZU6zxhWUsYxIqIw+wztMD9cCAZu0qgqZMMYdxPaxnHwEabPxTABn04BpHSxrTFBSALyhDBepxD9V0ML8GYC2JyFmCCrz2EbCNaFxB/IvZHFhIFrkIRjeqygRmwQwuWMISuSCU/yUINQRJBKIKOxhBMBRiiLv1iEc7MEYgwKEL0kFiFGRIRh6egQwvrYIEVxCH5GzgkTXYIQ26KF3pdMEKO7BCGrTcxChGgYQF8EAgVSLBNvIQj1VU4RmLs0OBsGEDGyzuGcAAnkJGoDwqAEMcVAhGMGYQjIVUoQriaELHKLUG62khe9vDxBvwkEWp0GQRNakJqq6RPp7cgX1GUY1RRIAuqNzKKc24C15uwgAuhIGQWCNWJYw1lmRZ4BKI6MdQ3hLRdiTAZwaSAg5MwYZFsMEULphDKRwgLnGRSwEI0I6B1OUuEbZLMvOyjAAE8IYlfGUPxqrELFr4QgXEEB8yTGBrLP+Aw9jsEATiaKMJePqbIX5kGkbckBKZ+AWOOQUXGJhNFanjBz/cAXwHsgYmHqCMLh7DiYc5j8zMGEgYxGcJDGBjAl4xNgVgAI5EmM1s3nMHa9xqGnnc44ICAIBjWKAI6nnCBw7xAqt5BGsSUGIiF9mAU+BgRH3RIAWa0hRWVPJFBZDRBN42C92KowruEAejeMGLXGyjCmN4RipD2Qkh8QgII+jBL+wQPVws0w4LaAIOriCCKxj3ClBgxAKcgQQpRAMXdjgvMs+LC/ai173IJJ0dYsAOKBTiCqBYBULoAIUVfAQbTnDCAq5bBWBUgVBUSGUngoCGFBgglIS6BRV8C47/jXxjK7VYhhYcgSkOdU8AcXBJQSu4iAnShAALVZ8FHHoUlb5vKKHwoEVtJQU5MECjHMBLRz/qP5GGRYAC2oUQRACraK3GBwoQhgOFgICZNnkDJhCFA3TaU90oAAdB/Uik4KiYAlRChDIgIVKVKgBMSIAJTEhhCzjgwg1U9TQyvCprDAZZ2dDGAl+wgBzCikEM9qWsH6FFD5CoVob99SNvlWIVa0QdLNx1KVvc6zIe4IWWmQcPZJxZIOGjKcQ+cmwiwMBGTgDZ6sixAHegxdHSkKDMNugYRfisBNzALh1YbUUnMUkJFMkVHMxBbCUqG9qckoootEgGTKhEFTP5Ni74/0EJcMhGIA7loxHg8xkKsQQlqABKh7hyCrFQgumUyQPomS4N4ABHDGIQgVSoOwZ2gPd63cteZla33rqQd/RiYANGkKEKwRhCHqCgiHWMYgWZGB04yJGQAyskCIQyQAra2U5LDEEc7kgDIV1SjGUAYcP+tIIKOhUAEO+HAAed4EFl8gFupK8nDh2Gi9si0RjL+CM0tjH+rKJj/p0hpCMV4AtUsAtBdEE1K42WDwqzlUesAAGL4MQiXLABaJhAA6UQRSmmrJs53OAUMl5XUd8jrzR4I6kAkA+ai9WCWfgLGtAYxpuxqpqCWeAQkZ2AwTBhAbD6hs8ZBI68GoCIHuCa0P9NtDUrPpDoCdRIindIkVPqYY0iOAIIy1CGX+fHHfSUkWZPgIHNljABNvr9N/39mRwY3592qcJWS0nD0phmGQDA+o9mLMAZ0nCraJwhibiWQC2u1Wvd/PA3CQi1UD/Cg2KXgQkwyqReHK+ENUQ7FypQQ/anIA4ySAIYCWE4FViJpBwY4xfq/twCxrD+N1k33vCeN77RK//qrpf+78VFfKfr7gWc393kBodfoAAD6wRCebiHy4AEzIJVWIU8eIVQCLPNc4mQcIQHwJTsUYEm2r2PaAY5OCibIp9ZwIA0UAUUeIEiWDFY8QEEMgoYewqbu7kau7Ec86hbwYUzCKBiCTr/FaABDDC6FRSYYdAAJ/iBrbgHOOCGa4AERHiBD5iABPABodC6nRoXBfA6sOOyopIBsmuQzVKBF/kKYlEz0dgAVCgFBMKqrCIECyiAoGmB2tg7PROrnaJDBwg8l6CB5GAbGcCYQrM18ZGDAZCiARDEASCELHIJVbAAIACCBwACv7I1jQCES/M89xgaIFCBHCA9TwuiBEC9E1C9xkuYDiCEVLuVOGCQVGyaSLCGRrCGOFCFWKSFE4AE6JA8aXgBFykBtumBWggVHNCZh/mL5JsfSOiBFnm+GNGL6JMDiaGFQMiFEciB7Mu+XEAGSRiC7zseQsmFYOARNTCGb1o/9Vu//3Icg+jBt/aqt3lrL3pDL1yot3bMv2SiN10gR3M0R0GpggM8niAwgE5Sg2DYhmFwAFFAipqbpFp4mg37uAwcjw18IHGQIJuaoG0ZwRJ8OWhwn6FIIJp7PZvDubzIiwmowa24wQACuhKIAgtAAQooinagIblgha2IAApAABxAgAFAAAZwAauTlqwTF924QuWLCi5LhAI4ygL4ALIzu/EAACDYxTP7ikRwAyWQAikQhARIQxlqC1BjwzacjSewgDjkxJ0CPBf8iFpIojJYArYsg+VAPI74hmmQBmuABFWgRUSAhGaABFy4FUUknAdwhGUQAGJaikkULJqRgdCbAivYRP8S6QJxgYeyiUFFo6LqIITKEqo1iL0F0SwGAYTQjINrAIRsQB9VsLDXg4Mz2MXW7MVQQQBf2xkNSr5biYBjPLYyyIUWoAreoorGEw5FjEYrUAMV6JERCIJtgIAhcLCH+z5g6MYpCIRYqIJAwEdzjAH1mrfttL/ufEd5S6/t5IHEuc5ybILwO7Ag4IUMiEY1OIQ5MEiDTAAigkGF9DgNwxQgEI8AgEga+8CZOhVCgINUSLE70MhnGYdoOQq01DinwDmN4iguGICSdIr+0RcdHCAVQIEbKAq4EJhxGAZXeISt8AcK4IQKYgPRUABZ2MihkLIueAUrtEXbNErHOISlLKH/LhQAINBDGdCXOzgDJQgDCoBCrEqNdhCBNXSP/njDsbSAAeApOty6KxC8PNzFMmCbtwSBL9iFWpjRNZCCOhBTJagDJVACHVACGpjJrUAEFcjPRhQAW1sDzruDSqSjWFhExyy9v+uLBmoAGquRGpmRDvgAzQSspkFUzbqEeqm9IlCBF7iDF4i86AgEXWQbFvDF8PGA2Rwb3SBGobpNJjg2ZOPNqrifqhgA6qOFNyAEFphGahwBSwgCYBgCZMgAA7AEA5AEgiiwYAgEX12cclQ/0Fmm/INHeJy/e4vHdSQdZIIvWpq/+oOT8ly/QWk4YGCUhJiBEbCCfUgHFhOFBNAE/xlrClooAvz8OP0UgLb6iAWQA5qwKZrihKwYUBO0gFiABrbw0JmblVAYpAaoKJtDAjlAgJ28Hy7IyTCIxELCQQD6n0pQSQt4ARzQ19OAyaOQLRURH05oIReAhg3IKQUlClEAPAqglI+MgDuYGv/wj0RYyo2Ag88UAGUoiec7s0qYADZIUWgohRnCqrdIAEIAAdwrAD8Qy70bgHSYwzp0gFfwgBN4Citdm11UgZV4A0NrAB1QPUIURUKsgxl1CSbMgRwAAi14gMI8jKS5NBbINDqCgXPVgg5QgDaKTHjo0xgU1LcRxMw8GlRE1EQVgGPABMEtAgtQgR4AAbq4EDhQgv/WbBFMDbFNDSuIEYEwONmmCNVRvYBSzYsBYIBUbYBVJYQZyD7iVAM+kNUgmFUqSAFeMIBaRQZG8D57IodfWCZaEjdWkD9WQFbw5E73YiZ444E2gQNmWsf1qi5aSrfxDEAMIAhCwdYMkISHQzA1YAFtKIp5uLouGFcYDN2y/bj8VKpGsBp3hdeZKhX9WQMCfQELcINVWEH3gQsFFQV/fcHD2AohoAAC2N/+5d8tANuNuMGQcliIFboo2AZ9jSi46IItmJ8IkAOa6hdowKme5ddxINk+PVlQ9YSVRUqkfNkGiFlEndmSiEpStSmqk4W38FnWENoIacOjfdIoLYXI3Cn/p5UfGoCBtWmRt7QAPPiCWrA1IQjEGTFiQiStWyE8TcG+s5VTta3TmYGBWYuFB4nbuRWryCzZjRCCGvnNGfGDDzCZC4mD8TDjpvGGwD2GV1MGw5UAFEiRxa1UY5MByOVADxibTq1cYXOJX7gDUT0z3MoLvEBVVd2FWIiFV1UDIhEl8JvVIEiBSKaCWm0Cd7gFDBiDNKiu6GEFVuCBY/1k3g1lYxVlUG4v0uEBalIm+1PWd9RdXQAHDHgn1k1AYKDeIDgUK6AEOhCFV9neTPDe0LUATCHm6xkP8nWJgT3fqGODjqrX9n1ffWVBBR0Gf92IgMVfjcAFaZCGOOCGNJCG/zSIAziY09lqgAHWQbAoAQlQAU8IhYqFlgUiIsSI4BSlOpAthSLj150KtmxugB+4AyJow4E+SuEQYZnFBE25mDPbgxYwhRaCBgfwWa6sIQxAgfSQATc4BBmwjSd9BRvWKZLFIA+IgI+IBhQwtjJ4kQC5M+YorS7O20AdAMFzCsIriUwEAjzoGI9Q2/XY4fX4gMX8Ajw4BjeouqX96AS4gfJQAq7NpMb7gEk9EEAYM8tYRTX+IkyAtRfAA0f7CDjIRSYoAbFmgUvwCGfA4wzqs99QAAp1ihP441FtaA6oCkLOyTOAg1p4A2OIhRFQg2lUHud8ZEc2gIdLATD4BdKZJf/dZWxXbiZk5V3vdEfeNV5khTfjtS7Kfuz1goPhJYgmGAPfGZQD7ATSHYEWkAVRwGD3aWBydQlasBlMSddjthpl1paHhjouqIM1YAV7dQMFiN9pHopq/tdgxoCCRViEHQAJxQA5PWefe1h1VgEVIATgVg0EcgtRiJ9bcVc24ISpQ4UKPgDTaIu4KAVZQD6b+wEsEGj/EOiCntPObBoyG1s9LIML6AAJUmGLHZgaIgQUwETckwEQuBcolbKCPPCmJemvRmlLej4f5tJasAOn0ARCpApma7zirmlBWyKy1em0tYZLQAEgxgMaQAQT1wE86LgCgAa/4NNXuIFoWIOmjj7/3RoAljuaRhCPqmYQNX41rYYQPJDqpdCBsR5rsb4El5ACD3gFPqPCKnRrdYnrCyDVXoHQAagDOPiFXeiBXCDdaTSGTijswrZlB0sIMp9kMhiD6bIu0illxsa327W3OKdsUs6/OHdzaJ1ze5s3VoCEVIivMfgTfgyCYPBrPtAGXy7vLnCsSWqKNs2B7CFmIKDtZJZICopX3eZt37ZuD12pF/tXbLYoTeCCiZQgmcBy+sGFKEBJHyuBHlCBQ9BK1UgNH1C6oGoKJBgANrtnE4g7pGsLrEtvGYME9h7oli0A6puXPaK9SDdh56sE/Y7oiU6gPLBoIPgsGCgAGBAPEBiA/yYP6Skc6aCCA5R2vnMvAwHpngCYcLMSBAu38bfxAwv5y8K7GK75AjlNg1oIALPYGESoBUTwBlrAAzdlcRfXYhjFARlvakG98AHAgCHXiEiwFx6PBB8vAq1+ECE/miIXa7I2649AAhFocrPsxLZe2J/5YzSr8ryQic/N8lrgcj748tPN1cGeODOfOGCQhCtwh2ftZDfv3fg7L91F3speR2ZCpsqWbOCFR2gVgkKQOH6sXjXghVVgsfdxgNqUlLBVgSWwgkjPAWMWAGQW+XetIPSd193ubWjudBaElmpOYj6+lUxAgBNlg4T6XEFQdejuMXVmZzl4BWkOQmpAxI8QAv8c0Nl+2YCeXKkEiothGIZhnyRIMIb2PvZkh9kEQVQAcNP0WMsLmAmqcwBa7+8kRQFYw+geGA8UMPBwj7KRLukGsIMX+PhRZQJ1fwMJP5B3r3GqkAOoVWJ7x5g3kNM48AYQWEyfnuKMBoFLOfgs5rNXwIEUEQQcqPGcxPGtgIMAUBnx2PGLPwa+4qsiUIacHvJ6KHddFFUYwAOPEAaS3ymdquG+qNzSUhcY4AMfZQKAyNWCAQMOBAkO8JTGF4hAuWKpGTHCkCUDQQxQsWjR0kUqwDpSGeJkgR1dPHSl0sVKFy5cPFixcokrJo+ZMmnO1BVjU7ieMUqysoNzqB1sdk7/8mgCQRIwKkGeBjGkJuKseT40YG1XygGFBg3WfPUa1isiFSxyLLFiRQsQAAEAgfUqRE5BNqZcmGIzQEkDXSheWPgw5+qBcQc0HNYgKtSZNA3qPRYr2esWBGwW2WVjcMAZsXEb4DqT60Kl0qRh9FAxQNThA+0O+xB1A47XuGs0WWazYQO0DSY0tHuN74CP2ONEbJn8WQohCh+efyD0vA63BmkiRQoQQIAATADeYCqCycKLARx0O/DR+gDxA10w0ABwDIgKGBIACPgyoIuDraJKicJfFx5A4pUdLzxRAhNlMNGgCjt88UYA0YR1TxhcDMDABBoiMIEciExGVg8KllBC/w4g0OZZHLWAAAMMMrwog4wwfKGMI0xAk0ACXfAHjwMO4PBIA4JwsaGRGn4gTYhrBHDMJAA8yV0kAhyjzDJWFqFMEXgoWVttKLBQIhMlyIBCXMKI8MpWW/3YhQkeKEGhV9OIpUMPMjCR4BN+EGSQQQxwEUYalzSUSys5SGQJL1SgYREVwThlUVMYUepRIU78ootKQm0KEw9C5RTTSqKCGpMzJ2kqlB24dGrSTKx8GpMdC1xRCBVOeeRUEMFMoQYfq1iF2DgaANhVZGB95hUtL5SwRFo5aKGFW418NhdBdrmA2V6g/RXYYMIWltg80JwRR4gN0ClZZZmxoRkHAwjimf9YoRVAmr2VlCBBDwgMo4F6ryHWBQXJeiWIZZzstttv7SD2WnGiaICccmJNs0YacGAMxxoax3Wddtsdo4IaOVixRA5h+nHeBumx1zJi8MAnHxBASPCCAAHo96N/DvxXyoAFNsAKgng2iGcOFmACQgCsiPUIOUVqyAACCAxABCIEr4FImGM2i6JkcMQRAAhuxFiADE/IEEsRRWhxwQY6OiDgjzicsgaRRxI0wQfVTQaHAMpMEjgA+EVySZVaalkEEHg4phwNLMigIBOx0BDXJiLIIkp/pfjsgAmhCJFiZF7R8EIP+koAQwcccLBIQQRxgQU3NBQq1QgzWNLJDI1GFYz/IRldFMRHGH0kCRWSFFLIGDyk8pKnr540KqeiwurSUSqZtGn0qm5/ykpjOIGM8Rp1FAQaI0wxAiV0zIPVVVeJ4opkBJMVRbPN5pCDGjfDJZYSciCAAabIyyI4sS1W/EUFgiGMYQDWjsVEoTrIOhdlDtauDZjCgJ3xklfoRRrT4EtfG/iXa2DzHnl5BQMHS9gGXgGc17yGPRATgSYm5pVmYCE60JEOIeqgJI9phztT0IJanMUCCRCBCxzgRBfUox72BCxmx8iSBIpwMzwM4BUm4Nx//hM3AnlFaE9oEBmZoAILvEFpjWuAPbDQoYNMoENEUMW5EHEHEpVhCV4TCxwA/xEJFMgokDIwmwyydCPf7KhHP/JAKtYQhjdyAVAdSlKI7CAAICxjGU+ahACmFB7EZcmKXRpLA2ggATGRCQUp0kQCMgeg/sTNBAqoQ7pIqQMWjPECTLhAC/zEOtgRAhAM6UEuZhCRTlDhdobQSEWCNzzhCS9XjhrCFaoQA5NcL1YzEQqsVNJNT3kzet/EJjg/xQN3XGEITZlU8CwShBmgbwS8kIVV1IMVUQzDFbWcoGRUEQUZLKFZz3JLHD7zPwbMgnWaWcQAhNAAO/wFBB9IAAPDdU9oeAIdFJzMukyxATa4gHXb8hJYcKEEN7jhCU+4QAFCeAcFzCNcADsADZeEAf8ObABhvIGGCxnWMoBFrIbzE0sECEGEAnQgER04RAcKcAbaAHE7AhhiEUuWg1xkiBMmIOFMBRafY2BCGRYoQgAigUUtco5YXfyZV1IRBbSV0YwW2AEILiEn0BDijQdhwAAIALTJ2BGPS3iBufjYCLG5QQaJNZvZ3GBIGbABbnJzABgfSZBZwJGSk0nDF1SwDEcsw0kAKNwnMRlKAaxRMog4peTKlKJMtLKLABKQAgTxGdugAAa6vABpetk61rGOC4RQhS92YIxYjMBXlAiGGmbQTmAYALrQvQh0gUepaN4KGVdoAg+QAiuYVO954s3eSpzXzZqYkwejIMMVmGJdj3T/xJ0SmUIsmDEM9RjGnj64gZCWJBZIRGFMeXRWDgj6GUHIYQITUGheBqCDh9IABXiYaEURAxxRQOMOdNyoWNalmw/rhS8cBI0OomA6yMGADyXogRsG0zIo0hQJIcIFBfKiU2hAIx0+CI5MDyAKH4jAoSQl6geS2oEjE2GpT7UOdoI4VS2QzGRLUIEbNsSAra4nMV6VzzHm84UANAIP4kiACXRWCmL5zAOn8AokeoC2MfLBQSCY8yXWiAtCRA12HSJAKs6lijsQTQZleEFq+4hYxQ4y0YW0UQm0mkgH+IiykHDkGzGLWb2NUiysAEEOgABawRVOcYpTBhC0JIDCToYG/yoIaORc6xXY8uzMZ/7R55RAvwa0CG28LUAvCwJcQFVBFbsAwUMk0gk+SKQVFzFAdJttieFJMyO5WufxJHEFMDghBM4AyqdYFStyYhMpR+mmpngADnCADxlDgO+kpBnNp6AhIlNoxSpig5XCaGBYrsCFDcWiih6ouAwlMhkmAlBQ/yXYPAzQDBv88GBcdIvC4DLMPTlxh1pwuMOW8agLPqoXIZOSFVHgbSVIs4cQFuAVrHkxYjwghRBFo8Y53Q0qeGrPEgZnHD5QAMjnRFRCdCDJSj2yU2nTx0YgfUpULVnJgHAHPwTwN/dumHso4AsuT6IIxzD4JeRAZjOrFUg8aP/rJSSMgi/MWQJnTCMedCGWU+B5r7DbWx0BPcYxRaGwYIHDYV+QWLQxVrFfwIQjYMABHbkpbouMQDTyamU4YiC1XpGGBSQwswc8wAtuwYPiZtZ5CwAA1ZKhhQpGsIQyMEiVr4aHLIg1DFnHLRS2Hp1YQFACXffWl78mQC120YNDSCT4EqFCRZgtieiKI/lVEAcwxLF8YACjCtD/SFOOXwhJ2OIWigCDDUZxTVRhr7zZQ0q4TwIOd7DXeB15JvnI15QZ9EoNvJjD1NuxY50jYM3+9QoPohBnri2BBBTcwRVMgm1IQrGOODwYK5SOChAARYELUImCC7gBDWRcBV2Qbrj/gF48mGTcQ9CMnMlVwsmtWCK0XrhAkQY4wdhNRircQLtwQm/gmCxwVcsYRigswEYV1ZEdmR8c2SFEgWNcB3ZkxyWpxREuARBEgRzMwiwsjIXBhmzUAn5w2dbFwSWIgwIkgJlpzlbgQCOtwQkA2tmczeSckQVYAB6YyweeAgXsFQdcmmYBlt0VTd55SR95Awr8HRk2Vo04whJwgAk8WqSFAiQ0Xp5lVuN8BitYgMnkgCM8wJMEAOepgKgBgeKo4bnQgjKgRYmUiR1QRhe4kub8yI/IHv2sge0xgQxcwBNUwkBwwdRIEgLcAA04RCwsgemNgBWMAB/wQvEhHyFoQgUs/4AzSEEEOIMzVEAFbIImbIE7UMANDEHyAUMh/EET3AI2hkATKAIZKEIILEB3jd95ddO5jQEF1MoQSJ+0QVv7tZPwdAL6TMU+pEP9YcWwUMNfURAPoEAUkEfp5YAKYMKpSQaCTcAAcEFCCZAcPJgulI4FEMBWTVwUcoIMWOD+aRwbIEzHaUsHhgVkiFwrjmDJ4UsPyIEoGAbLaQB/hYgL6oZO1ZwDCMdPtYbL6SDQ8SAPOpUQZkcQAUC0qEWUKSERTMAsJMCZCYtPyUZ8DE6XAYA3pAEtEIACKIAJwMNWKIbm4AANXII16IBuseIu5ckZpmGfeUUEEIDc5Q0WZJpY0P9AYsUZH8BAFGiUWEhDdrzAB6SUGwSeGwzeHxrljpQZf7yCAuhABFAAQgKKJHHBDehjSQ0bHrzB4AjA5hWBCtBH56nAF1wDCq1BLRRB/ngiCHTJFnQBgAxDPGyDAsSD5pyiZ6oiK5KGDIDANVwDN+DmNQACIBRDFbhB8PHi7XQCs6UAdB0fBvxANOBCNDxCc0bDOzzCO7xDM1SAMOgBPdSAK7iCE1xjNoaALWxjE4TALfwBGTgBGYTDGJzKScTAAnQDGbDDeVIAUzAf801fNLkj+VjC+fTKDDBDTFmYTw2LB/zAuXwGD5xBLMBALJRICbCAMpzagRHBAPgB1BSEHJz/AIS9gANKJAomhihwghugQAN8IIep0AV1HEg52LmE5BPUy0iWQBQMQHG0RwrqU4hAAg7oBm/s1AnCUAm13MtRUAR8gA8eWQv8YGOkASB8jFSpgBWQTBEBwQscgoLNAVIShrDgACJwBxUKgDfAgSoQADRUZZm9kiiAKAhIiO3x1gWEpRmBAF3hQS3EgWOgZZ/8koZggeQ1wDfUwoamRmoEgjV4BWQwqQCoQAEoaqKZDY0Q3hJwgSCaQJmVmQME2RrEAR58wYYCBgoAwsUQzC9EwRF1GhA8wNZ1FmbOTCUCwRcQ6oipAgDQxxHBwAu4XQNgQBe0Jh3sQy5wAR24phDQ/w8cMEuD6NIrIgAXYAgC4ECy4gAR5MLt5CIvWkEn8AKzYSv0VUEFfENzvsM0RGcznIMekGu5lmsScGcIbKN3Zh82uut3lucfKMK8yqsT2AAFhMMKUIC+rsAgRKMr4ADzSZs7Do8xRcSvzEM7UFxrDGiG+hdYpIIn7FaDlAgQRKhYCAIR+KCCAQoHYOhXNCARmAA+gAtiqIcDcEEPmMkFnqhOYRAnKOC5uFUrkhxpsAAIIABhsIc9icLAhMgJ6OgGaMNuzKATuUxNRsBG/UCRdoAPGukhnAEgNEJP3gx3POkRqoUWJKqVImW+fSgOgEAcxAEgiG0ccMMapAIFuAAqfP8dz/CMLHDCXAGACoQlb+3BKp4RXUUmHgSAEIgDQbjOnwxAHYiOZ5yAG4jlGPXAhq3BNGTDdqjAISjqohbAE/gl4eXABAhi4hEmz0kBAEVS6FKNX4UIDQBaieSPFjiCAOyCCqhdJWKmBLhqWHwGOlQmAGDCeGRiA6yArr4CFyQCJbQANMSDA4AOWJSoV0RDsZaBSPrWIiwRA3DCLDADL+AiPM0AL/JBCvBCChhAcWKrOGxBSzzCKTSDudKDuZZrDdTACnynun4nu7KrumYju/6BE6yA+uqvHrgCGUDfdWnEdAWBREQEJaxCv0Dha+hcKDQDCtHeKUgsb+EJ6k2BAPT/z1dkrB/4wUFCDRFkqB2E7FbhF5AqRoiCwK1NxonuqMfFbEuOnGySZAnEggvQKHsAjANgwLnoABfsaG/wxsoZLYx5gMOeC5EOQNP6AZK2ABHUgTcEkVRZLZQiodY+gYIpAIBgKVYMAyeoQJNqhzWsQRtyAipoIX/4DOdwcXjcCc2GpQyQJSZACHj0AJ+8juB6QorUUgP8QizIpkqxgDeART2sAS1Y7eQaMtn8pRVMgI5MqufETQJowgmkZSTBDqBQQJd8hhhGTh5Bi8UWgQSwgOu67mUWwYaRkjUAwAMAQf6wgAV05hr07iuEwiFQQifkAi+kgywLad+8QJg0LxPw/5q7DNASMUMLzAA8NcsMLEEwWEIKODMweK/3Rlc4SIF0jiu5pu/+YucPJIE7wK93vmu7buO6Zp8t2GsF7C/6uoI4BHD7CTAB484cDENrONAC7/JtiUXEtilvOcjFYrDGdoCCcSwBZOg3hOwr0HNr7BiIusEZoLBnYMDCbaQLcAIbyMEuS8bMiiXJlYAbKICHDocPdAE9nAsSWAYL4ZgCuE4ATQ0BYIEmaIIOFOiQfsART0DTdsASN/ETVy2iHiHJdHIVTwDbJp4JdIEChMI24EAUyEdTb10Yu6ELUOWk7gwXZwku7bMuuTEaWsCcfQcmPF2f+BpfYYE3EKBY/IIbtP/iLj3BHeCBBGVqZfZAUyWCIRfA5TpCDrQAIw/mI2/BCfxtHcMOBZilZIghXDloDkzBMVgAC9iHBGhBFVXRq04GKj/AMozMElhAYVFAF6wCF+QCJYh2LjBDOoQCEUuGNPSymACzbzEcM2gDLyDbMWPvDFBC90Lz9+p2cUoCEjTD+V5ncGfzdWInPfgDLlRABMTAGIhnOcdvc49zOTcBO1BzEgy3/tLDIOCAdLUzd0cFAfuiPDMswwKZjBWqWECGV0BwvewBP/OBCqhhXETDFhCAHMgBhQ7AACAAAbzcN/jChhLBK9hfj10YJzyBQ2fcGqjwBqQoG4gDamvaC+/zHpT/QAHMQUIPhwZ0gTCESD0IAicsQscR7be0jHpkuA+cttISwE1PwAbj9B18TNU6qRQDNVtU2QTMASzJlijIQigwdZcdA5QEQBjnFQKEAttW6o/ErTIoAwu0QpuytQxwNRrtACaAxx0sGANALxsUBBfEAiZ8QS0U7h7v0pPrkjJcQhyoQgDsAgB8wVwT3eSmzV9qwV6TGaX6NWAfxC8ZxAfclVicAC5RLP5MggW8SABKgOVNNil5hWUvAxBogR6ZyyMggTgMAS+IdqbzglJf5GQITUAxSPO69nmwARfwAfayQPbOQCdE827r9jSjs3AHtzAIQ/vSg3SCK6WfSvM4AxmA/4E4g6d4Cvst2AIYsEMm+EMDVMAgmIF2ZoIwVMA66EF2Ml+zcbd3x1tytQIXzAFrlCxsBJkDTxAreMJo7EErJMIePMFmFtY0RIMqIEK8y7s3III18NtnAgYRyOS3qweIFkAgFC4FYQBmbKTQWjQRL+IZ5FKbUvghmEAJ7az9iQBGF+oWVPTMbQAqDMbN7SxsbAMIgKkDo2WLs3hAdwALcMd2qHwUV5XJKEMPtACObw6xYIUGzAMXy0doddmQn8IHTM3aIh5/OIBVN/lKZTUMqABgzFWVg0csLNh5/JaGyIAy7IAA1CXpqPU+P8EU7IIAvMEXQMgXsIAfJBlSTS5eW/+BnTeygCQABnwunkKvQWBAWzbACehW0TCByTB2ID12ohcBLZzLNQjAZTvCKmOCuXwDBYiAH1hCptdyLhwCF4xoiOjCCwRUCaAeLykUB2gDaNN2CdD2bTtzq0ezdFGAMCRBrTO7GfSDE5jBCqxAEmDDI+AC7UfDMvLAKXTXApiBIvRBsL9vc5MnGHzjCvxAc9K6M/CEK5hBONgAGYzP8R0fs3k3cyUXJezDlY43fgGZUJESZIBFSF5ALjR+K1CCCuwCAeJCFeA0fiMkASQtvquAHLgQuEBRbHDCvwf8uQw8QLBxsYGgQDknGiRU2IBVlAtPLkS8sKeEn1cHNBzAp7H/nQ8RERYmXLOFEyeC0DagmuNjY7sDL1+O84HgBR50a1jFkbZmTYMfBCYMCDqhQ4sOMAAICKBUQFMBKqwsiTpVWY8JExTIElVKQ1evnCwAmHTsGIBjAdacIjRgwCIXoRSYMNHFAVhlyli0kigRhgoLf3e8wbQDkxsuHDiY4sCGAYcJMDC9EeCrUYAAuyxA3COxBJAdAN6ALvLmjp8OpzsUUO2mCCZHWlokSCDXgQkHXboQoiGHwazGixojwAAnZIMTMC4wSc6kjIRJFtwUkCGjhAQVEorUUtgzYRwBy7w8eKDmS5wG9iis4kWJPftOlFrlEregAfeE0l5IYFGiTAkm/y04mIUDbfaJZYYZSjjwwE5SaNBBBw1IYQhkVmHECSfICGcMZ3iIoUMeKkDilEceWYPECirw5xQeWIzBjHAW6CaEGUNoosYQwADDxhAykYJEXJJIkUUekMDABjKuQKYQSYChwgBgnjQgiGDUiIoXZhQo5YBhDhgHI4w0EEGT4rZrAJconqiElxlyKIGSEXaJo6c1cMHAD6NMG6CDCT5ApL5aXrCAC1l88OFLQw0VZYMCoiCuPjLrw8CtgQjihI2DykyIlTMe2usCFiYoxQcvXRpHAx88SEUkhR7BwNIN2CBIJUMPcCmmLn0YwgJMdrnsi10iIS4CoITyYwJjj2pqqf9lm5piKqmWyEEZFfzwYw4HSuFKFA2G0UAUsMhapqyz0sKALQQWQQUV2eQCCxO8JvJUBhUCtWAHwgQrQMDFOOAEsQnuiAw00CJTQTOJZJhi1ze+AGEHEO4gyrTUUntCmWUcsaKDOWabiy7cCHihAwYa6xcxBrCIprgT3EhuuRKWwESCAg55wg0YYJDAOu1WracB77yYZJkHtADAPPRC4cWS9ih5LxdKchmCHOK4SyWKJUrgrwwmKpllFm144WOGVmYQ+0BLJHRwiAaHuIIEdv4YJYYYfpk7Ah5+SMXDGFJBooJ3SAzcmXV+GDIGcHiwAYy5F+jjRltCsKWPMeYGURj/f+B4RIpMIoAkFR4QB4fuMZpwwu0hJJHEACqoHIGFfbDU8taMuupiC0gVsiOKFloZwYoRyngzzjlZoQBZPQcw9gNIGrinFhCiIIQQAj7AQBBBKMABAQTkkKOSKMzDvT4KFhGIIFg3EAehhXrChVOI4t2DCU5eEWXbjF7SwINTQkoDBSLYECsXoAQVJvBBRlxiqy5pYAAWUEZgLPAFyWQjDbtBwAS4cBVkwUBZTHHKFHIArahISwW8mEAoHCCKFG7LfqLYhgXCRZazwIEViKCBDnD4ghd44g5YuMMdBIOXVmxmMxGRgQXqda83EOYJ+zKFKRjjmIAJRjBfGIzBJLIZ/z54JjKYAAEILBCxq3TAD4moGBCU8ZpEzCEuc5nLK14hjh6MrGScCA4W0lAcHcRCIkx4AhNKoIwXFCA10smZBF5wCe7YxzuTENoDHCEA86whHCJYD9Pes4emyacKeayP1bDGH/90jRlciIWBxEY2PlgiA2lb2xAKcQUN1S0GEajl3GJQuL0NyW+Ae0Q9HhGNH6yjGSz63Od4EA52dGNIC1jAJhZwONDx4HMRyAQk3hENfwhDRP4wnN46JLox4OAKhQCGIUYwgxFQggPQSEAePIADV9xgnhQgAAaEYJ9HKQQOGCDECJbgu3QmAgZvCN8aUmE8iSFrAoRQ1RpUAQIVcP9iGD7gEqIKdYBSLKoH4cPdGiTlApNU6lIgWZWmOBUviRTABXMQgQfiSQ0c4IACW2BFQnzWgGJEwQ/oi1VKVvKSBHZpgeLYQRECk1RePcUPDJiAU69CFDd00ClNsUAInyUtZSRiAKF4RSlSWIphtJALO4ghWdBygg/IgQjnQsAAFTAHBIQGL08oYkSe0Jd6WQAEg9lBLvbFBn5xYgABw1cXd4DFvfBhCjuQ4Bv4agEYRJWMp1ENGl9TiTnMQS5y6YIJZMGFOZIMMYpZxCwIAQiewIG1DdBBy/YCSCDMrJDTYcEdXkCDRSrEO8eYhBfCI8kGfIMCeWBGCp7GNPZokg//vFDfJ6OwH1FybR+UENt1DxSMFGQgA0Po7oSuQLlb2tKWuKzcLlmEBCT4I3CPmIY/1lGBIU2TB6MIATtsIE0WiU4XMRiDjG6AgQUIoxnTwEU0KrAJXRpuSIVj0Si2sY1YjEANfODCKtLRFZjk7wAOoACkvhGGKvRABQCdwe+YwIsSxEkhpyAAQ/e0JyzcFKISRUBFaQcTUzmAAQW4wzXEN77yCXADlhKHSffJkCgU4AK5UKlmcdwOU2WkFDeohSriEAc46CIAPWjB+VyAipQYUIFC7ZIoxOHApC5xiZigVoAYwAWo+mGqVa0qCKG1hGgpowiJ8AMqXuGAsG7Fftsw/+sxxCWuAMChGeZiS1sWEQpUxHUAAgCAMkoQr0pwxgJ+sRcI3rBEwCKGE09ETAtYMBhVOzaxENk0kxnLash2erIYrJZpVKMCIGRMBkQgwmmI8AECDPsOMBjZUzkAHA5wgRB4KIYvbrANDMQBBbBlckQCKYFEtEA1BchrzlCgz+4IwJHA9YJw7RGOPGyDH0NYmnLfE5FYiOMZushGD7JWAuq0Yj0swK7YcsGL7g58CHmYzy8WEAHy3tK8uywcJIi0XhLZg0TvQFEMVhAOG9jADGRwghls8IcryA1xrFgBDlYwhmgeLpdJ8NEa7PCDJBTzQy0C5y5DcAVxpLMT2njFAf+/RDsNdGEFxYHDM3LRgxwAVKBWmAElVAwCT6blxUQ5lsQ8cdMGoAMFFkDAtryU41N1ocd3UMVJjU4+NpgkVlCUA5IXsikmXzsilDBBV8bRDqE7gAgNCzUeQu1lbWjjfGOmFf6I6gNRHGIHD1yiEndQjUDwggMki+qxkGJnp1xVz53PARCOUYAWQMM22Bq0A3BwsWUkeoYnoMCjIR1mBShADpbGBAvi5eRKPKEE9PrLXyKzg0PMYhFQNBkH/NADTOyKMITptKcuwAd7DWbWKpBBBjMosdSoII1WaAEbTZCAz362Lnc4duVN0RgusGYHI+guF7YxhAI4eTObLoEF5mj/lNrKgAXhzqlC0kAAfAu4HkC4HkHdVmEV2C0FLOE9KOHdWgE+OkE+jAHfAKkEWmEfyAZBFKQVWIm7vGsIjoAEwsEZEi6anKGWIiAFbekHzKtDKgcJLucR3qEGHwEXKkATYsCbdmluusEM2IEMQqBFOIRvvKlFeCACkgAJogEXHuEUhGETUsGbFmyXdKG/RkHngmEEeGEONAyBMMIHuuDDFCIVMKAKjKHERkCgAkoNIpASSgAEPOonjOV4isITpCEhAAEzvk7DvCQmNIDHfOzskiwkokHtYoXt2ODIyKQhnIzJNm0PWiDDgC7HEqAAdsBe7OWoYoELAugkxmzDRFED/14hF47qXlDxXpRhBPyg8ioPqibADZJC8wQAzzovWkDPDXrK9LKF0EJL9S4GE45BAOAgAl7v0RhgETghzFCh9gTg9pQjfj6l0/7ii0JtBxJhXxAjQJBP+ZoPsbDormKNzf5CBWCACwREg4ziELgvYzSrjbogAV5hLkSrA2bhqRgg/QLEDSJjBPaBFwAS/rQhEZzMyWSgCIytjA7hA9ygB84gtxxlIYDmt35LuN7BFfIgSfgBGfiBH5TGAdtDk1ohPmahEgwE6vggnVigAwWOu7grC4aABMhgAWjgBBUul8ar4XZwlypgHdgLG0jkG3DhFDQhAn7gFPYGmTzE5qYJmf/ma0j8QRMqABe+4ZcqIBOc4RR48EOWMpxCYEmMYQZ4IR3mwQ+/xAFugDhUgQL+KaDWUA1858TW8GlyAQakTiEi4AYuD1n8oA7ycA0AAQ+KoA/DLug6rCRjgWfETSEOsXyWcRlNgRPerhHPgP6yqAVkoTAzQibmIBYeKBM/E7ACSKRO4u5eglaIihQ/YAocDxXbLAp4QbDgDINicRY1zxZvEfRgoAC4IAEETRS6gNBQDxOKYPWWoQiO4RLgQAoIAPYQoC2W0QUIoCkAgAWiMSJ2jwV8rxqv6AkOIRHMKBF4oVoSIdW+sfnCsY9U4BQzsdMMwze4gAsGQP8kYNesQLP/OEv85kL8EMDY7tEVGyMWH8gfG4QXUoAX9mEf+GEWEuEJYoFeigA5ZzEAGiEN0mAN7kEkWAsQBCBoHGkSBAAQGuAi82AVkOEIkAEZIAAC+IEBQVKTRDIC96EF1kSdFGQGOqElsyADdpRHSaAJFkAKEs4ZVpAH/CEGWJDhGq5wKoDAaNAGb1AYpCApt3JIECecnhIqP+QHotAJScQfukFIqIlvepAHnAFJgKETRmAI6EDxoGAzD0AUbiAQCGDC3HIGlsBG4XINDYEZOqASSgAFPKkB8nIvj2UA6kBl1iAO8AAE+lDsDsBQHIALLsANamExF+IRENGnSiokMjQVPGHT/0Q1ImZhGPIOUcIQGnogFVFxDVmgB3DGDWTgEKDhSzasVEzADRqLVe+lCHhKsBYBMeJzAgoAAGyzqnYghPRshKbAWCehAEwArIQTrLiAOI/zOJNzOZvz0Z5zEdBFOi1DAEbAP5iAiKbR0xxmMKYgClTA0xIrEzFhV9uM1dLTyfhADZKqPV8ABkrGN8aoA3pg1xzhHWVj/GwDAczvHklL/dxAGaZgCnhhFgDyHwESIJlBG7jgDnSRC6qFCBKBId0gCgDBQtMADizUGjqUIs/NPHDhBkoUGcSgDVJURTvyI9sjPlqhE5rLElLSRnnOJXk0aLPgCEABSE0wAoZ0BXNy4f9wCQYH7AcmzgmpskmrkMGG5Jjmqyu7kkU2YR186b2iEAY3QW64skOycAikxBhyYRXmAQrKsiznwJTiMp2cLk9/J09ngJX2IRfqUlDxUi+zb4z6UmV+Bg++AAG4QjMPYB66YBW4oBIsNchwgQIWI1YEYjEmcyF8ZlMqYQ9E1XO1oVv07ktMBQG4j1VLiBda4E5uzQ8UAOgUiHYS4A5ck1WrIjaN7xUHoFiPdfOw6hZVYBLcoAXYoPRUCKwEDQcAIEKZtwiUkznPZQC6dRG89QPCtU2Y4DqfgAWQ6PcsoDV6AB0Rgw1MjQN4wRuRal4Vq8mSA18frxzdYGHnLPmAQAv/7pON2GU/HQBhOyCDFpYDWgAGkOqv9uFAD/QfDRggZ2EVBi8+q6UDGrQHvCHL4iANpCEOUDZoNFi4TuEGZAMCjkBmV3SE+QECMoAXniaToG5NDMRng2C7XHJHZTgLQGEmTRDhjtYmbSlJy8sZusGZZq7igBJwuFQKytZDtpIHldJIPySJeQAShCEJcAFw3gFIkqBwwsEJRmFLb8kGriAFxAEY+CAYtmEe5iEeOCERDiSd0ilP29hGmysF9mEbULgSZOAuE0IKcEDOnuoqWgBR54RRBzMzaacj4mEbQiEBHvcJaCDIfuAG+kUZJZkTxEEKPJUhQvUCKqEAOpcSoOGA/zIK70ShgXhVDWLTBSx3A0wBFRyAqEQRI2Z3V3lVGX7V+BjDqYqVFmvxdz1vEqKgA4pXWktBhQSNC5b3OJmXGKGXWweAAdoCAbAgEiLhKZagDGQge5OjB7pXE5FKAiYgkhVDsNigA1TAr5oPstJTi9z3Xv7iBTqxMUjGXx+jfrWgAPBX/GaDP83Pf7+5nyEj8iYvA7gAGbYBgQUOQSs2PgePGXiBCHwsAKwBECRaojNYZQUgWH5BDmQjD1K0hFdURUEaAuJvaRDUuvhgA0fAA1sJaGc4C1KABEYO4YQ0BqIpaVlQ4WgpBjbBBpqgG3oEF4b4BmkwRG6ubJnSKWuuQ/+WmGtnsIpxQRhqIAJwJAREp+FWwAnQNgWmRCx5YcLw1Gdt9HdGIBYMoUFO+Aj2oUFzQQZQICKl4Ab42Kk41g/OwFHS4BLwAAFkwVs0YB5kYRv4lrMmYA8YuThyag2mAbHXQBpKloYsOA1YYRoSQrI3tzI1WZP3oAMUwCtk4lRUqANkeRPf7HxG6lpq5bRd4lR8QAFWlVdb1Q/IV7AUY9kKABOS4rYtTQA47xaXIHhHIBGK9zdNzwFeQXmB4LiZ93kJ4Dm7tZmbeQI8oRGmWQVyAEGwmQm0ea+YL3wr1wVyNxHWs3aXLxz3YDOYAF8HgxpVwDBKxjHu8TFUoEoKIK7/CtYE4EEe+3NP+pi0UG3VYoEZ5AEUBDwBC9pAEZpG1yMgeSERRiAQLroRskG6U1aDJ4FCaUAcZCMdTBQZRPijIQCkOXIVMoASDMEQTnqMGWS7YPglhVYE88AGEO4EbHLGkTYn5yZHwmEF9AAXnJCKnbAZNMEFj7iJsTQJGYxMyxa+kuAUDswJhUFGwCAcdNK/CgEZIiQFDCAlczQl2VhB0glHLWEfvEtCsoAfDmHT1rqtFUIHcEBAGmMWMsgPlIA77voLuCAdZEEW0kEcUmksTWAAIiLcxEcK7EkOCOAGDn3YCMGSFyJDWaEOILESNu37DugLa+cDXJtaUnkDUGIO/2TBVk87I4ZhFVrbtXcgEGAbigIIMWahA2zbWHM7KZIVoIAXAFQAuKP19G4DAZa3eZdBudnCmZ9T2AcguiujCLQAa65bmz0NMPDvMGIbioIVvM2Z+jrN1eJlHNkZiQzDD7hAdTuWF55AAuz3AlSiYPP5FfqTCK6Cn53ZPJUoF7YhAQUcFFZhwLchA8Th2yuWPcRmDcfaGAjBGB6U+8oBuJSiEXZBHGYvAQR8G1L0w0e4DT58FfhBHDqhE3J2JMsaBF1SxWVYaK+AEdwhSBdAxpE2AqQg5Rdu4bIQDEJAGHicBoX6CZOAQ5gYCVnEH47JcyCOTEUn6MsUCUbhB+yAx//9IQnCAQzyq7xwaQG8WBKwHMvR6eksoctnIBgMwQAETsUHjo45ucnuOCKRoM25kQEQYHXnPCHSIADsfA60IRdY4MtbYVDmwA/mT9DZRyHqoYMjczGMjxMIgHl6Bg4Q4Q5EVdIl0YDwblS8JQHcwHbbD9oTsdNbObVJl1tCIbxNnRWjXTZngQiKwFhxuymAQFlvMQee4xCCOYWG+xWMGQiKQPZlHw/SQAfkgLmlV3q3ZwDOIMsiARO0IIS2hvfaVbvvhbsDKLYXIxeYL32dTwUiYu6ibz39KlDYtV68iDjJYhLouQTcCd3j0QQQwA3YnTadigGSbzA+U1A0PA9IoN7/QSEPQIEOQIEECPpA2aMVggEgZsxQQ1DNlIMEBfLhE8tYLl6cOClYRWcVhCsWSUDQuIrfrFyUQnbKFczSPnlDMqRcqTJDhiwvs8DMQ2bMggVSFkRY4EynzwgRYjiLETRGCHY2kuB6hwvXo6dNK2yKwOMHj6tYecSI0e2PIkVG/ohV5FURGLNmwXxaq1atok9g2LH7M3Qr0a2ZGA1JwTdFBirBRgTjRaUTL14ZUuxN7FIlsiG5KlXaU0kGCjgNMgvhwoBDZwYIJgxAsaYBHDi7PuQaMcLKDNczeM0ZNmdCpVwgMGeul7nBmt+Qbphiw8kFGxemOBGAtEZaHHSNauF5/yGj0gXJkme90jBOg4YD3ocp6FHkzQ7zO3aM4MJmQ3sX0DbMkXWgXX3w9+dxUjElvf//gfjBBgdsmOICBwh2oAwAAuAhAIMM7pBDCUtUOMISKkzyRQFsmFCKA6KUIooDDnSBAABAFJFiinikoYMcAwyAgIwTMCDjAGfEEYc3mAChhhUllMBECRJY8IIFSFqQHgtcEDjccAjmogIm5+1A5RsWqPDEdVzy0d8bIOyA5AsfcMEZZxNw4QcXBbAgQQ5PQDNHAgmYUGedCLhBxAR81lijHz1QeeUOU2xDBygkIAoKKHksumiiJJDADzO8WMLHDKwVZNCmjhzk6RQEjTCDIf8PHWYqL5RYQgmqIVHSiSUZHJGFPDKxlNJLuMIEEzIkhLMAEjrg9NMCQu0E1F1BxdWNP/7gwoOz2DjjTDfh2OAVGWC0tRYpyJDyiRHghvuJt0asFS64456rLilkEBvDL0XFQMZjfvFlQArBCIQYY37ZOsQ221wn2RO5yJBbb5sxsMhnDEzghw5rpDHGM8YQqkZros7ABzPxiDKHH3vk8gJm9zRQDxx2lJZZcJwQZxxybCzXgCq7gICeCiVMhl0lHDjgnQ/deSdKKCrsUI1/VPbAhYHtcbKBfPR9J/UB3Q2z339Y7xAFLxzMwsYszCA4ix8qAGD2gwKkLeGFFVaYwyT/ALjBQQIkitLFhw68gsAXRRRhgYpFtPjijKEhYPiNZ6SxIwAPaKFFhTKwoIKRSf49RSyzMBARG4twguAHSu5QRJViasmldXyoYeUOIBz5ghsMzILgImJz4YYEFcZ5p53w1LlIAXv6IRqfDPgRxdGDTmHIKvE42uiizzOa6CokIAMBM1nwAkwwgY3g6aaghh+qGgK10kpIqqqK6vqUAJMBP0eIcYSsut7aUq4xZUFCHu7ctMAvPonBsCIwFKAEZQHsSMZYssUOc31LXRAs1wPVlS5yncuCESyXLZB1l1FcARmKqVdiLCGQGTTGfi4ZQiHEkYvInM4yummAJhCgMAQx/6BhXCAEIYwRiO9djA8GsEQwcpGOedDGD9eJgjQyswZa4AEFtUiDyU4wAA60zD0wk9ka0LELMYmpOhfIRQEkw4FS4Mc73ikFApShjPSYxzxKM4V7NgAf+ZhxHPeRWjtEgQD++Cd0YlKGCkbAgh4UspA9UEEUjIaJN5jtbDuQAIXatoS3AQAGc/tQiEZUor2tCHCCk4NobERKGd1ACYqLBAAm0bgcTKhIIBhTLAkVC85wrkCeY4AbLNDG9FCpdFsqwAWE+QTVXQlJKoAdgThgCit2rU0lKMMFoEGnO1WTEx9IxAQ6wCcupKkDPQDAG45mHgvEIhcUiZ6j1gkpjUCAH/9icIm9DBAEKhjCEJiagvc+NQLyaawVnegE+lKVKljJ453IEEMb5leIQuCKMY1xia5eMoQ8XGET/huWADcalI5uZRSMYEcG1fWHcIGlXGrx1kkv+AlG9IIUMIXpV9KyFna4xQhn0Qmy4BUCvSymLxmwBBoE0ol9pFAlhdjGFmhAiDAWIBfXecLBfCMIGnaNDcyg1Gr62U+DBKMTQUwBJQyxDVmIQgMJ8MMYoxCHzKDjDXiwmS8AQYsXDIAZbGhPe5JDABpkQ0e+uJkMnsCEC2zpAtoohXfaMY52eMcBAygCJqrxhjfuAAZNyisdnzYHM+pRahoQBRf8CMj/9MANqC3/gBsKoBrUTgkTXxBn2gTwBSC4MgdayAF/4MYCBsyhbg74UBdMpCIgfDKUM2rYImiEgFOmcpUPcIQacsCCHFgglrFEkt/cwBlOPGlAXIgF1tCTJcPuIYyG5Q+VspvMzgyIc81kQAGiKU1q0ql3vUsAJwpwiG1OoAXdJMKUxkm6WBSAEtpo3qGg57x2RgoZyKjVECRhgApTmAoGAAYwqBCEehqCCmgojCUsYQDE7AtgEEgxhK2HjDaIARnzk8lDbzVRmcikEHkAw68yaixi+fguBYxBOBjxwJPCZS1wOcsfQhCCbqxDWtjggR1iMAZbNNCkzogWGMD1h08oYgF2eAQu/7CBi62sg1pmsIFOC7iTX5DhCouRJ2M6IZCSyMMl28BBBNbwCzdEhmBhlGoM3bENvFaKDyVgDWv0WRJeBLHCKUADMGbTBbQisQAw8AUc0lALm4UJBJiwgNIIpNe8siERKgATekSnAhjwgQmEvcA00ehYxo5IDsqY7OrSgzlSb9aOZzyjBiCLJGUoqbRag4jslsmMWbTgtSD4wi4A8AUBWGBCS2DBEihkSQlw4bfBDXeJtlEEFQDub8gdgI0MR7hTblqVk5jEMoDwOHN/AQTYVdIUYKc5J3GCAeHdQS93naUtQfW8Tyia37BkJGNklkCdQ9B8mVBfE3Rhd3TaLxH80P+BAQhvAFxANSZG/gYqWeAJYywAM+iQh/2t8+WIqh4E5ifPFACjwgagcIVvznNI+yVWR4AwBKyXYhUPfehtgHCM6ydRGg9BJnfOAjLy0AQk3CQnPd4JR3e6ABskI1vWcjKUyfwOMT+i7E+BSlOccdKSKmId33jEPXjQZSz74+yPwEbemXWKGiShGQQUIAAjMAonXEGEck7MpWbQCl7w4xmKy0afAQ1V6zwjEBiogjgOkYuF8KEVJQwGGixx8wo7Guf2ZF6INDCHFgyzFSoQgC8EECbS7aAHE3BmXg/EBgF/wT/mKTcYrSOZ2SwWjWj9ACaUQVnk7UCZLpMjsKcGWsj//jFrWhMQlAr0NbIV4d5fcGRsi4BtbVNIAnBTwQTAPSK8vWIbb5AAEF7gNyB8IQ6DUzcN2Y0AObxAcY0wWw8CN7CFCfiWJH7zBDe0CIswIM3EBXdgNP8xBcamJZSXXn9zXWPiBgjgJAXSTBwwcbAGDRaXABdnJwngAkRwCBznMN0kcuNUWYTCB1yyKnTAci+nTpGyETAmE4pxLziXczincznHFxJ1BElXdEXnTkbXYvGzdBQlUfhjYxkAClfQDTsmLFlHLENBLEEhLU5gA89CZs3SLHrnFGRndk+hdzFQd+hiC2coZrgQDkZGF49wd2WIC/7AA5mQBEPRDWTgBCJg/wZYGA55ABOJF1GWEgx8UCoPkQiH0QK8IImsYj6fxwfBEAvB0ApUYAlGGEIpAIShmAKWYAhckA4gUgri0QFh1AojMDqs4x/9cXtcMAubYyDDcQhFgzXCZx0tVAkdYALeETShhVZuAAAk10hUAn1O8x6dFWyg9QpyUAT9cWxY0wPaZxwb4ExkU1k2I34AUASStG3kaElFMAB00wUkIlxdwAlfIAHiWAT09wWAoARykFwycjjNhUpxEAlps0rLsAxasCC0lW/lVgAI4jmc4zkD0APIlh5ZwgdbgnJ7kHDncWxGwoENaEUbGYJCUlgbYHEleE2HwIId4AfCIzyHYAGTUP8NzrcDNFh5BJNgcwBzjhIpD7ZQDpUYoSiEFhaERdgXMhF0SqgR7kR0SKd09JMrNDaFWVAIoOAEWYh1AfRjX3gX3eAEK+Aseph3d+iVZXd3afcU7xAOWwYuXxEDTlF2TiFkn2ALYGADznCHeliXe5gEmbATghgOH+UEZkkCEBVRWfB0KUAFmDgDjGg+rXCJaMAHhuCYfBBQlsALiiEPlsmUibEXo3gvaCAbIxIiwwANrJgLTCAB2AeRuKd7BoIgqJY1vRhVldAC6UBr3XFWocACjYSMyrgDCAlxyMFZivUdeDSMGvAKRHAQYrJq/tEDvFAgMJMcY1M0YIJvsMU32Eb/JNwGN0XgB791N3dTIibACSAgAeTpN98XB/aYXDQ0AItgOHKgA89lNpNwDPO2DAyCB/cWS+WWCwkJJf/GBT2ANFijAq/2BDLwanxQNPeGJK3DgczUgBHnkYe1Aa/QBSWIgipYAB1wktwkPAVgAZSFjEczSNnGAiXAAiiKTvGwCouyYI8Sc1cwdGLgg0MAhEJIYTg6ivUiEwrVBm1QlEuYYj+qlIWwlDWWK7OSAfJwBHQgCTeBBDnRE1uodQe0FSHgBJvAA9iAh3TJpXfnFGnHdmhxFmNwD0xRdnr3Ds5Apt+ADe+Ah3q4pf5QAeGAFD62AKMQAmYgAuzwQSnRL0c6/5gpQJmORqiDyhdGZZnMIA/bsKRZID9HYJkyNpiZyRfaYwkK8ArBJQqcCg2keQFMMAID50UWAAS0aIstMxwNqItYoyQqAEbDFJuyQJxCowEeECgxqIwWwJ++aSB25APUh0YJQACmSqqyuAOBIAfcp1ecEJ0QqWqOJI4UMq1LIAHHAADKwJ0kso7D9QruSJ7yN4/oeY/smY/L1X86AAf9CCHxJm+TIAABAABxBSZfYAHKRDv4qiYBumrkZYGGZVgJWo3Z9QJ30CS000wDEoKDJWsUOlwnmHEr2AFEsKEDcJIfCjfIKE4Eeli5gHJPcAcWMAQ36HI6uINKN5iaKQmjSP+EOpcCKpsCg5kFSIiUG6GETbhQkDqpKxGoSQoBeRACGUWVPbZRXngXZmAGMeCmXVmGZvelZ1eX2PANUvsN97AUaTpmT/sUeUiGelgVPBAOrkAsK2AGTuAKTTAK/9MHjJAPT9e2geqUtEIrhfCUS7qkMTY/shKpRhpRiiEO4rAN6aCpIAIi+7UlidaqyXmqnAChnsMBrJo1OANVHVsJs2BW3HG5nIoAIOpIkzVOFnAIneFdzmlH3kE1aHRWCfABvWQBypkegUAEi/te0Ek2EIlv9GoBkhQk2bYEI3Ctx3AI3Wk3eBOeIAAD5Dl/KvAFjaAEN9KeoAEaCEAE6RoH8Sr/n6sENwEQAGmzC+GHCSpwCLPjTLRDu/+hagU3kYaVcMfWOg3ageEbXwUgA7J2ARtQIsM1kqggB4cgsRvagh+asdUAADtgOv8aaJITBUQ0D4fSKCWbYksHiip7LxHssqEYZzzKYinGhEwIAUPqYvLjUPVTY7NiY4VAAldgE0E7QEVbtBVgBuGwpXlnl1/ptFCBd3GYhlyqd3DKtWWopWN7F8QyBtRiA05QxEOWB0PwdFMYE3ErszaWt3grP5D6hPMzxfQzqS7BC6Ggqd8pCq8gCi7QsRfAByPgH2FybHBUi7HbOckhJa36Bq8qudfBAcPQHcTIqQNgAZMlTpTlvaDL/0xWNBxsMAdnRYzEKAIfgDW15x+v64BQ4hnk+wL4Fkv1mrsnSiG4uUrAWyLruK0eULzkqQLzuLzkulzPKyPSqzjxOoDXC6+RkL27gJ+hBr419G+xQ77PepEbW8DqO53XRbCcga8csDDyJb8MW6H3e3EJgAoDMLHOzHF+oIvXSm1UssuytiV8wAJG8gEIYCjxsMCM8ihH2YNJbC8ULMGQ9rKJMZQzm8E1684cjHQvBoUx65QwMbc08aQZJUDGIgXG4gwRIAVb4Q5Y+ix3F5YznNAHbcN456VPS2ZkeIc84A9vOodhu1FI0A0rMApom1EL0ASM0FD27MR5S9J4e9JVjP+3MCY/MIa3NpYFirEKr8DFnBxchQuqZWx7WJIeStNvsXtDH+qaODO/16ENq1erH0IEmwsALulIKkAEC6h7i9BZaGTHl6sAbgCLOu26iYAgzeQ5zUq+Gohv9TohuovJyvAgT6AAJSK8JOKtFgADPZBIL6ACIGAN6al/52o4BACf1Ash1hsAkfDK2kttAGABXV3LN8QAvLCLofNG5zu/T9DLv9w6BdsZVqQwQA0D88sG4lahdIIKH/AFpP0F1fl9DsIgseW9sUAwHMsE2kwmN8QG0BAP38xOMcfBNMcvm9kXoiiUQJeENWuUS2g9HTw/klpjSqwrWbANGTB1Tuo/Uur/E9NNpRtlA2bgDGO2tArd3WaItV663UyLh1uKDUKGtD62hXiaCSvQBOEQAjaQBxHG3E2M0lGMtwuVUAvlYvutUPPc0jFWCBAQuJysjuqoqfsFa3wQKFVCXjytxuKLIE+AbKwbxxdwXokADUd9uaXwCodgNCXnSAH8uqDxb6I71YplyMW4CsbwSw3+HyqQCJ5DO41bPLsoyZIcbRYwAjIQJCaabQQZC9BQ03jjAKFgJKR9CZcQAJeA1+RKODeCAARwAqoMIWgDAAHQCI3wyv8IAN+72AwTctIJfKtjTq3wr0+QoLX7y3egbp7x5jf0ATCAchwiuHmjzAowAB/AWh+w/1p+/gJXLk4WIJGGVQAeG9tl8hkR8Qq3rSg7OHT0E0Kaac4S3Bc/V6RCF6TEXXQ/6qNUrLP1/NK0kgVXwAjugMI3Ud0/MRSsHgGbYAZb+QO4cApLy90OfetdmusU7Q9yyus2EA6sTrRatwCbEALu0A3uwNF/IAJw9tJDKbNPKMXR/oT8/WLWDmNJl9/xsw3zswrbIAIkYuD2W6G/M1ihKigyaFm4V0P4ekNuYDNkDsclIGtQ1QGEHJwaUArjUAoJEAu6hglmM+J+AHA35DmmgOKXa9UiwuKDUllv9AZf8L3vKzZinW+V3OOXjKIEeQfaMFw17QAmEAovgOP3hgc0UP8LgnADhKOPMtJXaaALq2zlWA4IW07YaYPYYL4IXIAAXLCS6X4e3zjoEjmRvYxvOF6wNKTZi/0BJRBMnEDTw0UnCiBfK5gIGrq/oDNbZsPa6OuxDvk6hgPWnbMNr6DAkAIKQqqTNGrpbM8XP8WjCjXccr/BPurpeJs/Tjm38oBjn9DRKTylq74CTuAMezjeMbzQuH7rtV6G/vAD/iBkrsDP6T0sC1ABCzAGo2ADinC2jEACL6230z7FMJZQpO/fbcAP/N1iqK90o88PhBAFbL2tBt4FM40AT9D0C95IDv/zSpM5wzzM7g7vloUl835YLXDvxSgipaAAdxDiuQnwPSD/DoazgJqDAJ01DoVcjKIwDqFwB7p/HrtfcjH+bwdL8UXDvpUtaogGAz7OAgTZAy7g8bMf8i9wCKh1BzAgygFQBzACEAMQCCSIgAANOHECABDQkKGASHHiNIoUKUBDC4e4cGHAkQsCLodAgHizo+TJNxb4tLrwpCUfFSYtgJhp4Y5ABggYMOCw0Q0Llxc4vXJQtEuXBAkUMCBCpECiQx0OEXEDoqEAhtUsxGLp0iWfHhZeuNm4cxGDs1wIDaFD5woJuMjaIDuSJcuQDCn07uW7d8gQu0eOIEMGAQKJw4kRQ2jDGAJhwYLtZshC2bJdu4WyFMrjZMFn0J8jLBgdg/Tp/wgRYpix4Q/Xa388YvOI0cwftkeu/eXmvds3rt+3/Q2Xjc1MuBimYzhTjvrzJjLJnCj6wy5ZskKa6x6RJ1jMke/hB4uhi4y8mLnp27Thl54fXTEQUpS8s6qLg/v3X3Ux8YqLmxKekGEETN4o8A0ETdqhhwF24omDRUByQ8E3SJKJhZYuuKCFOURxYJxSQBSllFACeeOLNwBIMcUe/ChrJwQinKMUUUTRwEZRxulCFBfuONAkBIP8IiOzHuRgFj9UQHCmF0aiaQQZSoiyBBZYUIahFzjh7yj8+Fulh0MKKAAGGCSQ4JI65BgIgQnWHACHg+AAZKGrHoooDkAoukgAC/+I4GICBzcKiaSTKEwpFiaeULSVWGL6YqQmbRqAIxhhfAKoPS6Y5RVRuojnKBOU4qSpqZ6Kyo0v9mwIkx1iUdSrC2QIa6yPHNxpozsseMMYbehYZZUrIODnu7sywCuFIfriK1kjKCtkLsMQWywxw6pdDzzJMAPssizkyYI7wfIIB4nQPpPCueWUY26MfhhRxIZwVthkBREOaIcYYsZx5QfgcDmlX90A7hc3bHDhAZcKFFnBtNFKc86ZChYAgx0bQhgDiW6cYOfbb7vLQrzv4ENvvDbQa0+u9QprrDDCIFjFmF2qAeEOBfJzYL+jEvDvCSkHLPDABBHs4UUOeAJJBgv/gwRhSBgyvGCCDkOkkUYHPFASaBUBiIWXWiuFusYcbZxaFE56qAbIINMmktKiO0qyJCZpoqkHPkqoG4Yqi2DIAgReMaELov5WyhMiPihAhjJfQFOOAQoiaAACLoHjGjodaiiiNPDUMwAQDpmgTUA/4qIAQoNWcCsmWlKUD12LgJQmTybtKKeOuLg0KC5MwE+U/XSeY1SnwgwzkTtSvQorC6J8VVFZxbrjRdo3MmZJBHMBZZXH2sj22GT16h5Z8I21y7zGHos2WGpZTk+wQuqq7H1uMcuChCu6WYBc0M49t2HSnCkthiaw4w8DVEQeRHADfSTwAPkaRyZeU7CC+eYR/+8AWBLMYIbrsOM4n4mBahbAsA+e5lzhEKD9hHC/EDCCH+DqTmQEU57xkA89KVtPDVf2GMKAQhwr2sXManYUwAWxP+KAgZRYIIGfGUiJQpsApRwkoaQJyQIY8sosTOChEY2oFA5AANp2sSKtuahBOuHIAObggCyObUdXMFva3AiAjMzCibeSgwpAsIPXjcQCEqhb3ahkJYwgwAR/091+TKCAOzilAG6AwR16gIc0NQ4HjoOT5Ob0kOM1Ig2Zk0gjAsA5IjQOJLUbAOnciCAUoU51fGjUDh4FgibNbABtIiNI/gOUlnAhAfjpUlISALwCCC+Yd8DDRfYERzIJ6FUyiP8CLO/QRNqRkQuxAEE1glQNAERhG6sAxQonk4UU5CVZ4wRfssT3rSOsJ1qKSZ/55AIZ912GMt/kWCHod7FyLUB/p3HGaUyzAI39gQx5uMENzGEOeCTDBt3IRDjCAa9whGAFDOVgDLBhGhtcxwYrCEcykJOuEDqsn/9cATvI0I0x3A8J5HICCdrnnciITHsyVGcNzXfDatFhCIH4IoIE8AY3KOBvR8EZUhIwABgsoQQlGEHW3Figoc2RAU10Q9CkWAKnMYBTaOTqzQZgEhR98adfIIQ4/tSRUQ5AAWjMT6ewuI0esOqUSvtAWXRCx5i8IRCw5KsFesCzWMBABlUCAkP/QCDIBGxJcAogXDA/8IE7RAEPnmDcmxr3phsMgAKIkJOqrhIATXJyIhRBwQf84IcJNGgj4vgASVCEIDy8YRco2AEM3PAEGCgqFrp6FAqc1APGgUS4k/oAC1z1BF3yEohIcYEcCie8DxyCmMYUwEIsUEQZyOAJiYJBLG8iEI9M9T9LC5KKVMCCEWyNH6vgB14oE85yxjcvgRlMY8onrcMUxjAqWx933ret93ULM4XIAB3IkNJynesEznFYBFZwBTCIAAGDOGg8yBAC0iRHwzGgzS8+Mwp3rIACZngXBpPBDkWYwQnHCQcFIroCDIQgE5oAzRiiU7EaLyClIQjWS11o/x4gn8eGjlGZ+dDnK5AQwbUrisUP4RHExCZFHCVYQpWQuKLY/lRokxKuR/6zAxUh6It4mOKrLsCGV5RiR2t2gAnkENZdxDbMpv3TWSfFhTnMwW9+K4osTJAOTtzBmqgMUmx7WNc2gZdNRLBjhfiqx/TCIBZGZEFh+YRY/vjNqB9wbuE+AINHhsGyksxsZj+AiDTM6bMNCQAg4JA5TgIiEqWVQwdmORAu+IEQYXVjbEEQCxm44basnMkrY0nZO7OJC8QFiqImsEub5cwFHSBCqQoQ3RdU95PV5RMLShDYV7GgSS9oUaLZpOyq8Nq8eDuiCqbQg1xsYxuFwAtg4CvOcP8CBjCDKfJb2Dmt7MkFW0eYZ4AD7K3t5IEMOg7Nucy1gAWD0DRmgEIoCmBQeIAhBJvoYMdV83GPdzw5H1QNczw4mhqPYRSjkKgNyBAPRtjAHSkl10qFgATo5OGlMJwpemY4ZJa5kwSgoEMohksAknxRRUHdz5N7Z1Q/lCAHVWoqQ3ahoi9+kUGCQiuuZPtGEAClFU8oADSIwlZeJoAAKOL1T3eQC17cWiAIQIBzCXB3IsgBB4y7gRw+0IO0fZHXeABBXRW9kQHwQkkpcdILfPvXbwu2ShbYGwE84IFQYF7zCPAEtRXZSDxgobKXbRzjNttZbhszAHHY5CYlkicUuKH/Kae9rDhQdSLcq+i1LAi2DGLxe96CwLcjicLol73sAbihB9p9AtSWixSkhKLWBSCA4R6bbW98cttvqBKZGHkpx4OgRZMiyLInUBWsr0gF7FZBDqaAiQAQAgFXuAKwrjDvYxkrL+cUDLQO42+A06/seQ/wkJ/4mSf3QYY8aAL8aTh9gjh/CqEmUIeDGgB4ECB3IDmR2zANU43kADmTU5fmaI7R6CfQaAIyMAN3IJeUuphNwABGoAtsKQ8hQw+UcQycaotVoDscsCVxEAkeeoMmIyQoS4o5kAMWqLIcUAEAYAiGeIOf0ro32Yhzm6U7gMIgGTO/egJXKbum45KjUIAP/9C9FQmSQ/CDxvmTgRAInekSnOmSshGzFUER3QMBNxClO1s2RnsDwnMS4QMBFQC2SYsSGKA8PmGAUEnEpBCBOeA0ahMTNyAmLBi1zOK7Gzg11GM1bYsDOHi11ruGRog9vCMCPxCHAZADYvo6Q+PDHroD3+u9QuTDP/St4rus42sc5dMuN/CDOdgSUIm+WjuE6ru2Asi2T7KIi/iCHmABvEGcWBC3kWgRHFi2SeICszqEF4gttnuDQLQyCVCBIhCAD1iEy/MATvAAbQiF+tsGZNiGYhkC7UinwgBAxfA3a2GMkpFBegqw7ZAHzSCBBWS4BnzAz+inhkECMqDAg0oGMv+whZQKuZKDyJALQXRxjn26H4ysuU3YBB1DAhfcBCeIwcHgt5l6p5qqlvX6FdYSB1v6CPIDwjF7A0JQgMQSHKOaAwVAQglotzoRADwQgKt7g/FTw/K7gzhjRcETP2UiAgV4w+UKBZjhoV0AShAIpTQkv0lJrOXipVfwjx7gNaXjwxMBAUK4xVt8mzcIP1jyrRcQxOwqgUI0LF0SgaQwKrokgFrrgGCKxNAjPcaRg77zO85SNeoKAMx5NU+UCB3wBEL4gLuTA3EoxV3bhS84SqBEkR1gxp8AtlgkPN+iRas0RdL7O9vaxZoZKugTAemTCkVygw94AcOMzWTsgZ3kPd7/6wG1jAKxEItHGwkUwYM424VurJIeiAkBIIBzPMfLQwBz9AACQIFdeIYqEAdx0K8i+zcARJ+bEhZ9rAsCw4wMQLh6IgFGmLmMdMD9gbgxoAYROKgEYIQ/cEjm+ECJBDn7jACTa7CQIsgFMMHQqLkFuDkBHQNJyIMrAI/zoAv2aBnCKAxu4oQdQhBPMCvyOz7Wki1tlEmafAURQAp4SAoFUABxOCIWUAEmPJ6fDErgqlCsvEIA2AUYfdEe6oHbegKmRM2j6NAeiUmg/KI+aRw0BNKsxFEgSgATGICvpMwgBE7Cu0Pyq8YB2EPPnEVAFEQpgUtDBIEBSAC6pEsQVQDR/5MDOTiEQ/iAXZtEHKhEMXWuG8CCwSzM6sKcNIgGT5QGzcm+bRsrpIRCGA3KsDMuSWskksADFPhMEIgCq2wcU0TDXHQDGeiAUIC+KPtQBTjFRKi+x3pNw6yIihAAZawSbzMu3aRFQmhM1/yAKngsN3iBF63M2Fo/ZlxGFbCA4ktHzOOEK+CEUNDVIRCHKviLI5i3zSiElkEf/DrWasFB7YkM+cGM7eCYuugMjjwhAM2fB5QCTRABYkggfVCoP3hI5tDAEGQO/8nP/tHPEuzPfIqYzwDQixmDMdgEIZBXHiOBkQQygUOGKwCF68kAXoiFSOwBkgCAHrDK1EI+1lpF4P8kgBANUaVo2FAQURL9xuO5iqvbhfFrnNS6rCuMLeD8TfFz1F2sS8Gpy0WIAhgFzhcFziigPTR82ayMMiAqWXEAvKNUuj4VADvUWKyMUgtAgQqpEENVAUYSRGY8US1VCl+iyxDFS1KpPizQAQoYNSK4AQKwWiLAAM5SCG0zpkhIAzhYA7Gl002igReIgh64gztwA0LIBUKQrOD0WBgVmjsIrMC6g0GFzkKFJbwcgEX12wH4O+OSASKAhqQwILsMhSglU1V1AxTYVE4NADyIAhXogWVM21FFgeL728hkHEIAAW2cW5tQ22WUAL+6AqVgGWRon+zQN/3Tt2/5Dmgx1uz/XIygkwvykAzNAM/AQCfu4AwzgNd82ieDBMltJYYDSIZ2YYdw6M+OE1eIxM/lkN5wBaHRuMj/xEiawzmcm1ch6IYrYARiHYyUXIVtEAdjMIa6fUVHtVllDCU0FE2/3TVWJDxPeCxMJQQM8ARPuIMPUD4JKE4VYLVPugSf/KniYxzOHQBPSJG4jbNDZaQCIIJJWkPMgpNA6FEHJlS/6gFP6AH1JQRj+IAh4FJJldQEqNmVDc7fTBEUiIVTHIAg9VsieAFZLNQpva7Iw5tCnMo3EAcRoEkvfVinJYK7uz4UwAMduAQ8uIRLQAREgAQohgTUUz3QAttOzOJXM1v+bUwC/5jgQ4gCAMAD4ATKMobRtCWTWHCkvC1U3zoDAjBFBY5hwQ2sQ/AAX0ospq1UI8ZUtn1cTq0IyTVR2mSBtLWjN+5bxonfwAXd4HzRrWABRzJkygsET8CBVRCBefPHywAwAEOn2ZUWuGCnauGv3GXWg3NW31XAJqA5jLRW/amAcBgHfMmXQRgEakDeA4AHMwgB+wmh522Y6o1A/uknh8vedlWpAZXXjRyFQqADuNiGISCEQFhZBFm/SLRbR0KQbAqlvwRcOSAE4BQrFCCAIOZSpW1YBSAC2ixOVk29hvDhF/jgDzaG/vWEZ2gmJo3bQwW3RcgDX7LLo8o2VqxMAJgZQv9Y2zsghP5NWzmoS5mNsjlgZwwNTjMOSmMQ08ta5Br+IuFzY9/aikB9xlj8KTlwWKZVilDASwLoYzN9Ab2bpFO0WqzVWjlBRu0DLS1GzC0+27Q9VQL4XKAc6l0IgLiNgjtgN0OuaEL1zENYU6gOZ7RV20PYhlC4aqteTg/YOwIo0/8lhMelCIqwCDwwUUK23CYhVDiW41Nc0889Y+CcmbS1XN08znNEgG3QBlC4AmSAR9iFXcvQDvLQL2S13Zvqr2yhp2cVA44hTwxDsFcuyNAwg3vRh3zR5QOAAgyLgRd0BVcwA1eQlw+aTxEMV/5BuXxKZhbsSBcUAk3YSDIQXwj/ON+Urd9ASGpJMy5HUtkoOIQY/kvnMga4BoFcQGlfokkFCIUwrlwT/Unt47afAoFAOFsLmG7rHliLhuBAzC0EQOchblqrsGg8eNGMlgM/yDsxzTtdEmLv5tJ1ttky9gWi/qk70OhvFoeOJlQcduOZkTS4ZEYL8OGTVoAgLvCrbmkEx9QXIAAckOmCutq7qwNUk7XYtIhIcLWwFduwfTVEQIEXmGf/ja6qsFgBkO9duAQYRVvLjQXLBYE4S2IYX3Cozru8+wC0baRDYE5yJMdtuDwXiNIj/mo8iASxbgRP4hMVeAEViAK0dTz9xsuozjuhPvGp7KEPdiRHYlXk9ADm/+RBD6g/uhiCbaAMeOSW/hNAxRhl/LKWmXKhZn1WcDmCQthr4QXQgTzmFRiHBbLsAzgAauC4CFQOlXuoC+oHVxgFDtrPdD1m0LDzAEWCZY5XIRiFgbrXVSCBIYCZqXyBOzCGHmBxFo+CyhQAwvGDqA7ufSZUhmVv5FZN5S7ObxT1nC5goLwD/BZTU4dMOfAEMn7g2IqCNS6ARVDaRVRpQghOFDdjsjz1NVUr9i521fy7HfD1uH2D+hYH+z7Fjp6t2drvmWHGpJZkJQFKho3YEI3YA+/jIyaEBW/w0sNaCiAACb/pCjdMDBfbNdjwNECEPmRytf2ABpbcA55KX2BStP/9YMsVWDKGcRrYW0N9eHJT21xAgOSu+HNXXDkI8j8mciM38kjQ2d2k3GY68UIdxYw/+SkvcaAUSrrugSjIxi3Hga1GgB58k2dQAgwQ82ClN/h5IX44HxK4dFI2jJVJj1PmmN7VDt/NAp1z5Tu/1tAIBzKwAURPT3RVjW5wBSeIl6xXMSdYMVfw5U3An34yQXdl7Y7cBEkfBU1wZjqQR2R4D2T4lVUQB2r29DV2JLgVgN5m9kPg9aJeeAK46gIn8Is/hOKkXBX4gq7dNsmNAnFg6TXF7zOYyiY+8SZOS4lfhHNu9czzhKsz8QBg4mWn8TVtCrUKhc5P51ev6Iu+6An/RW+oJoAX+AJCna2mfjxJnus7UAEfHnx0r/jMuzviV3AGT9MBeHACoAAKqAMqljVB5lRX03B853DP/PAu5nXt84UAEP0UjwKEZ3IXxwMawH0PJwdPsGf19wQsiIJAQOoe+ACKR3fVTG6MD/JSHfKON3JvAAgBFkAMfKEiCggUeGig+EBAzsOIcgiBwLPLYgBfIHpw5BjlBQgCnDzgIIkABw45OLBcagSoUTFft8Jx2YZs25EsR45cQQbhCgkIJIYKLQrhKLI2SnfuzFIoC1SoR3A2PVLoSh4zSIQsQNJ1AdiwYKWEjbCALFlnC8yaXRDCRj8z4brVqAGrLt66sGC5/3Jlxgw1M/2cDHZCBgwZMjZshAvXpMmWEBiaVFksIg+ypJl9cv4JahUoLoeMGQsUaNcuAVEOySHSGiJETxbx+BKAgsCqUAoUiNCt24OHDz0OqniBJwDy5JcC4IlChIA4ca8JEDB+6WJtX5dQRLnTg4CH3btF7A7lIcrFXdct2iYE2zV8IgNChSJvv3zwHiBS196VEeMunlAnTkQEVocHHijQQMMuCqGwUQ/eedfDC28I8AYB9GmooQfUUXcIAR8QcgYBKN0wgBw3UEcIBYJAAkccjUQyI42AwAHHGjniuAYciODxBR4v6PDCGZ68gJwAASTpX2oXBRIFlD1AqdAlNP9UuQtDFHjooUNYvGDBR4QMcYUH5nHowQ0QhSgiFihEImMj18gYAAhfgADClxYoeB0KhGxJwHNEUCQAkxmhICWiH6Egzkg4nITDiTfc4EktaQASB6YxIreLBYTwUtMqV3xGwiokACUUUFdAwNlNyBxxk1VTFVKIVcjw89MqHohDTiDkXEHBGEh4JVZYZIFFw1nJqhXDApu44oQIZgyShF52WXsXttfute0KfDlxxTaFhFvIZsj0tCq6mZGrWRubpYuuUKCBKw4Wu6wGG6APfXCGAL4wtx0hZPamwG/meUBIFAdZYJwAkSTnDXJ4kJgvvgfO5p8vCYKQcBWc0EcwwfT/4YCCv9kFkFqf1OGr5nzh+RZyKJy4gR4e/WaUUb+2eUIIzz0T8syI6i2oEIMMRdmDJxxZgDIFZJpZJnAEaBnimiSaOICk1H3wgRLXwNgI2G++GceOazSQI4+IXIKgQi+8UAcKATh8s8kXnQFlFFJGQfJ6NCzU0JYgUmfkCwnfMQBwwBkMnJpr8oyH2C4BYs3Jdr5R0C7aMYTFn2oOyt/JG+EtZSAo3ICABwg8OkBKBCjRSKaZNoKkALUnKfcuWNwwBCceX5EbuB5sA+42xQ+xDQLbjPk7mR407wRJFGyxhRIUOBHCVl+BNewCFYilljObNGEGYa6s0E226Wu7rV3b/7o/yArUhINCIAQcvw00v6+Sxxx57L8KIwBYqlSRqoClAg0C53AFbQyAAKfBg4ACFRECIIw219kOBZ4mAqglDmHFWVjNkiNCiVHnOQR6zoFw5i//oKBwLwDPx+gDtRuQjFDMwVnKKJYvCshBcWWSIX0QcIe9lexkOcsOodbjoAYlaCELYQiWuJO3COWtQrapgg8X1yEKfICLIhpRiSCFohtoaWtdgxEg0qhG2OXobG5cQxxo8S88bAcFSkCBNxrhjbkVEUFPisKTiEQlof2NEA45JAUJ4IlAFC4KxhBH4iLJOKptDQt3gBzY0qgpBL3hDXdKyHKqhAU/balLKLgO3f/sdTcwmWZRqHMUSlIkKSV4Iw2xS6PDkmS75EBQRCIiQBXEMaILFrGFhKvDDXBADUitoAaaEEYFkFABaApDGDXAgRk2sYkFjIGbX/GKV9bhDldQgx1OkJZe3LeXa7GTfepU5yAGQQ0MKOQZVdiSSsxDJqc5jxMUQIEO6NcgFJAMBbsonJQ8gbfTaKcODsmXh4bpn5r1SZIcBA7C3IanmtFIbh4l0UNLGKL93NBfxzmolBj1tMUR4BJ9ZI4AdMC5P2lNDs2D2tNwMMQ3vLSYAtJaRAlwBjr6ragMkljekkohC+2CEBYlSYe2RgGfWQ1SkiIjBTCAAR1wIw2piMOlLoX/qTS00WxmTYM1vBHK7eBBB5icEXKKeIlLMPIMgTiDILWjOZf2iUV+YpFDCPcRT/SwJIb1APQg4pCehQGTL7nU7Gp2kQdV5BK1WFsYDsnFRGIBBHRjDgrwircXlC6ZTkCJiVQkVFrELlNIUpIII3GJMxACC1VYLAXrgKUFra0WNKheOFyBgUxUoALNcMZxm3GOZhi3AnqgBz1qMAgRhGMTSLAuWJKQCb+wox/9cEU4atCtd7qzndTCC3lhMQj17kWecLuEJxxyTwok86nAWQkqjyPXANBvoVGwK2pmi0igEkIJN1sODT4AVYuiJKMgeUFqaARXh5GIlB6a6inX9lmU/0ahh09FAAVsVkR/5ZBLISIEJO3rgQFIqYYjvtku6pDIAf+TqFXyBQ18kTEluPAjH8GYU1F339R5IKtYwAAhMIAFLJBIHFelLwWyutWuYkqsmUoDjt54tjhCLADLoSMKavGSsH12rnjCK5rpWCXf+pYGo5xqFfxKASOF9gUCOolJDIsDqRmSZ1h4xiXelEmwzu0ShEqQZQNw2Tr0eaqOfkbcSubSXdSVSC+4YzJRG0vVKsEacZCGLWXnsLnJ7U21QEEYwsAzEU31DAvCsW+x4IpMaGKaxXXGOXDdjF1LoRn0UO8K4BdPV4iAHeRzQndFID9YdGu9exnvO9lZgyTQY//X1q5AdNv3PmardxA3cPUlGE01Ld0AqiWhhrkxMFebLcdfCCZoC+NtndkS4rYUnCoBIO3SG9KAEHguyStJggPClQ6UEo7EHvm7as3yjGQlvWGDoFRfIScOB2H4rL9qEQDaUs1Pi8VCYT2A7sNCakrtfvgKzxDnGVOQEFSyEsx1TFfSuk2Q/MHCv82Ng6kmeclLPgN9ryqpKCeZqzACK9IvRVazNqDpPLoGxBCu1ox4o8ph07i7L5GQrROUNpethS/ATgNVI/kDRzZkHXSgA7wKSNOPQgnReY4FT1wij48ltAiV5K9iWAMRtaCtL/2KAUh/1iJotnRpNZ3MoVNACaz/jUMadGFLQEjYozNqxKnD4IklI5lnQ80xDS6LAgq4QxPrgGZxjbtc5OpBuvF8fTypQQ34kXP2ruj2enPPbfLWRQ962PUPmvEDZwS/+MqNbreaHezYD+KOEJSzQ0JO8tOqW9LWDwBDzhDa0IIgEPumLZzljAUDF7HfJ8m5YW+AkC846Dgd7WifRtnnL54S46GLgifqS3Jq3KAO9tf4C2DBVElVF9UWJJEcSSyT+mnffp2cxDhaAW6Ny80VzLGZL+zC4aEZSV0CzpEcalGAz4UBFtRBGAgCBTiZK2BVlGmV0YVa7GBZGznd2cDBS1gDwkldLVhDGkzeSxRDJGjcchDU/x29AP3MFZv5HY7VwZHJ3+CNoBCGFiFAiqZ9oNnV1p/VQaCBjUuAlR4VmpfVQi1gXi0ogQguoZI54c1gXR3dEbzdholIoZNFmQ7oIKhBHqbIiNhc3qXQAg2cQZFs3pKFgRL8Quj5ncbRAAa4gjCsQ+o1F3OtA7PB3rDJnjxRoiSy13qNl7ZRW3EBn/AJH/GBYvGFInO1HretFyXeUQAEAhOyiDhMoeJRwFzZ37tpn/YFAgicwVzNlvzxXL0RnrudDBagxDKhxNt9GxEmBEEFGo2QGQosWW3VFgiGgZV4WRqeTGjlH2oJHEoQgBD8XwAoAdDMH4vM3emgVjGiVnVoX/8oKZo1mpQS8MwAJllt1Z9lhZ5laUdd2ZEg0YCXhQEsolYVpBoWpFqqVU8cYlUXsWAdviDk7YgbOR0NNoI1UCRF/qDSVdmYFYOi1RER3tFpWBYtsBkhkiDnlSGTCaEOxKNVLZ4UGllBzh0W5tGgvQRcdVndWQMgqMIYiqBPYoCqwU1GxISi+cIdHSW8EcBVWRWUUYAQXEOoSd7kaaGgbSE69KES1IEg1IESCiIi0MBXgqFvoRoFJEEjnsM5VIBdSGLs9YMlLt8l6p6zTVsFIJczREAzREAoBh9eBl9y2eVxDR9zVQC1rED8uMIg1IE/iqOSNSYFSCEsykH12Z+/ZN//9mmfDhjhGSwhzyjZLcDN15VMFGbaFEoKXrXhKUkYnHgDqimhzxUkNWKdohGlL2QjaU4hBeiAOwajv5BhY9IjUHrCYwYk3NmRPV7Wbl6WDiBZ2clfm9xjLfhd6OljndmiQTEHQMJiMhECV4YBCXKlEmBAlI2nlE2PDkgDjNiSepINHDSde0rkmFlkRXoaltkhF0ZCMYAhai4jGPqdf9KAIBikQZKgEgyNHT2D0CWo2fmk5gkCIhSDFqrR5XkDxHhDGF5DHFwDIOjAVnqCd8Kmq7kjGGrHfhJU0KVgCpInCkBlHe6gpWghjF5KKjDESirBGXynDtTCCUQnctZmIGDA/wqcXuoJQzcIG1wOgne5gh6knikKWzwFG7PVAD0sqXIp1/BdqSjuGvHZpWAC5uolF2HO2gpQ4yr6JOc95uJJSktiABhe43IcIrzdkTLOojhCYyAyGT7uJoImkyvgQJ8unlChppUIWlWeWnd25RWGnaKB3W7ughLkn0u6JBaEnsYB4aKSYQhCo1Y+5p9K4eK1yQvMVTEsRzHk52zW5mty3pKF2dcVItidmnFaZ9xcgiCoaaTeACEIQoDqqq4KgXiOp3hqVRhsgRTY4Xru4I24p9lIJFipUbMCAgzCQaj1IEwUg4EG1CmFHSKowrbSAiIoQYB+p3cKIo22UBiQEbrSV/844OqAciUWhmEmpRGcSBiEYgqGnsBWiiuBUuqr6liJjt66pihWsSBUYopUvugaiVUaXEMtBJTaKQG4CoISRCci+GebkeUiThM9LF+wBRs5DQI9pOVZVsA5rEMSJF83mKUj5tqXAqbL/iXMeqmuLVcFZEKQrgAG0EAx6AAJMih9paCkAK2KqFst5GdM5Cej1qac0g9/9qTmDSi5imXRjt0NCK3VEsB+asflFSoNaOWhphoW5mNMJO1vQWqCpmBsSq3UYqqAiqCNBp3QkcHQhQFB5ZjRFu2Igh2qGeSfwSal/kJ0emstjOQTFpyCeJkSCF1L4irESqwgrORyBquUaVX/HWzBCbQoe95IWb3nDLZW7NwI6O7gYwFCLXjD0NQmDeRof6oC61asEGwlr3qtDgxN6pogeTYlBmwB7NbBGShB2EWoFlZk2FBkGrnoCXBoVu6uEOxopSItQc2ughCUeLrC7UrZCWCosdqhJjkr5F0DLZxA6qbuSgqCEGwrt4rlBdJAIFBAJgjDc4lXElDbCphPcaWl/TYi/nYiyaoec8Ws/74sAMNsXa6DYTaDeOkmCuxqdwoglKUrGbEp3t5tqcZEbQJUG37h65agBpNgIFAq0natA0MZ9f5T9EKRLwQvjP4WuEasVk5sBBdDNpSqjunAuf5surpO6UYw3tbC62ql/wYHqB01sMAqJQXAjQ6E3QSXagRvR3fuahiQQx2EXeDSgrdS8Vi2YUD54xhSB7oKLBYIAbiCsRJogg5sgVadce5Oj+UaK5bhCETKYNPdyA5mL6ZorhxP6+RcLEMsSHSyrh+rAiS8Lq+usCAoyIIwhO1Wr/Tw6iDTAC1YpBqpUUWmkacZ6/EqQY06LiYj7Q4fcurC269Wr1Zd71iB2hwjXWulATeoAi0A8vmC5QlsayqMJC14g7+iAJDSwzrQg3MlgfkIQ/+mnjPkL/7ebzAfM3J9Kf8ulxTMbP8mM5gO5skmwTmcrBD4lhKQw+5uAXmO8HiGARgaLS0o8YgyhAVDr/+O8TDsanMJSiy/giHVUgD1zjOUbRW2vlpLTLJLUORv1WjvrnA4Fy2ElmqV6AA5RBk9Y1X5egMtB7Q6lyA7b+VKynMDN2URQ5HGKfEEiyUK+DAJhqsgUGordysrj6XDWrAWK4HUuAIRY9UWqJ0QxLQOxPQWhEHupvH0aEImnADkuajmoo2WmRWPSCtRY9nSnc1Qn/I1WMOCgO8hD+4fpwLrzrQmiDH5YnIsH3J4Sm6wroAgxDJY08AJUDHxjm7CapJRpwEizDTkNu7yZgMtxPAHe/LQaFVW3TWQ5u4JcMNY9bQLOqSLXsM1tC4iRAAinIAqpIJUw7WF1uYvaEI4rID/NfVFEjBicw0zZtclMY9sWjLXMB8zzYL2Z+eaI152c3WiYVKTV1vr64KrJgQoBaxAbFfvFgxuMcT1ONOCNYxkmx2yIYvl+DKyruoAIsj1SAKoIgPr7NJ1GD6W5DC1ELS1GF/zI9cCXMs1GNJwclOAFCACFe+2bYPhGESscP9WKItygYbeQFsDGNYyLQOocPOqI9+2H0NCSS8I9BKULwDuqW235Z4AgAf4CbiDGavxFui0IGjC5apnG6PNskYkUsuxHf90hIOuRh63WK+Z+Uo1Oij2TMc0iMc0+B72V/oqGp9xi6idDhyv2nm3NaCD5KSRhoYVWCHrjUDCCSzAh4P4/wKcADrgNlzr6CGfwCWArxnj7OSmMSlDXlfN8XqO1Slva8WCL4DrgCqAw4+jQzZkwy/QgjvggAiQATX0BT1QUyNm9jDjr2Vv9v2iuWa7OZy/uWbX7zSFQyZIkzCsQG3X7hiDaxhkFZJz9RZ4N0MHeXsPLl0/9UiCsSaT7+MWd25HpwlyNbBuQfgeMuA2QjbE+E7SQHRHNyYrQUwPbiQ8sqljnqf/+QriNQYgNitfd6QzOiGDsXkDq61jQHpfwiPDcG7f9m2rcKOPsSOz8h+zLh8eMvTyccPermxHWRgYOyBLNSJoAoIfOK1V9fKa8g46uLJCuNm4MY+EO0QK9R1jiv+3/kJYorsqXINitzskqB0S6EC8f3os66iOlnGBT89NV7UURPe8e3cjwLhOYij2vuCOwEEqRIAOSIHa6Xh0n0A2qMJuB3lTC/nx6nuB47SlFzwbH6tP72Aq9B23HjaAX4MuxAHrbjkFmFM4mIENrED8VpOQbnYjMqLNs3nqiaxmd/b+eracD7POq/nJrgMj5vkW8CHkgrgmnPiJD7oqwHUj4HbUD65v/QKVizXV77iogzhYUvGPe8O0Mz0aZ8JXLkhYhqFOPnIa8eTCzy5MA9SWazpca3kj+B0N46xdn7HTvzpuW0M28LAYV7WoF6ivAnpeI3kYEHfo0QIgZIOWRzz/e/86xA4+xIKxi/vxYLMuOuCYU3syoud9oGPAV5+AFJC+6QsBtad+VWM7JLAxhcvggwu1gwN17CN1NEgrynOrKvyC7id2KujC77NCKjC8jp9FvPe4dxt2BJzAFmSCgatxVc+0FMS7DrRywBMvwfe1jesIK5B827P49W45busoiYP1CTh/8z9/8y85g7e/X6f1V4V860ZABERe5OmAGbCDIrR8eAFEpiQDBwoTtm5dhYQVGDZ0mBBiQyQOzzm0eNHZRY0Nha1YUUGPHmGZViBCpEMIEiEoNW3ZguFlTAzuMiFCd01Vtpy0GtGqZZIGohM0hp6oRUuVDpQohTQVElQn/zpV1hBpgokBK9aYmojWOiH0aKNsgADFIUtVx4m0a5WKFatTZ89aQsJclblFkCq9OXc2UjW3KdOVC04Ieak168s6OhDROAoIHbpsbnmqotFUiZDMThHRsqYqVWjR6IoSFRrUGi0dWVm/1HQiAuwTkE6cQIJE0yZNuFXeVpUGOJxoa9Y0KH7ceHLky4s3cL68ARw4ceKgi6MXkaoIqVTpSuWdW+gIUghLOSFFSlpIqrLH1iQok6b4W+RvQqIW/wm9gFRdG3utujiAG1A64tbwLgKhxksPNkDG4iubzn6p5RdahJIvvgzlE0QTRKgDZMA04BCRxBGlOxE4buLgDjRIRP+MwQl2bLBFERtWGGiTJOghaJ2DItqIoYiErGAiIBmq6MgKKkLSSIa6uVGhCoRJYoWvbEtPhwWQyCQTl7zsMpO8UsHJQak+S00VK70SShWflFpAByTijPMEz1SBDBBEDHOpSy9d0oQ2RCYMihayIDMLkGuEOo9RKYhqxJpGbhrrpr904PPLLboRAjQyJ1Olp5OWWknOBfTs0h0/XcJAEMaMunMqWP2yBp1aSh1VqeykCg2c0KYy6SsaTEPkMxpW9XIm+hKMAJJlI4gzpduQkGLaBVwMDg7iknOOW26he665bruVDjgBfU1lvVTiYCU8aVhJpTbz5EWPWfbYOyG3fIX/0ITfaRutbb9CrzkUHOqCE9HANd6FJJUIYosNtupw+sxekyKgxT1NkuBXN341EQIRdQUUsEQRozlxOHIH1CWNVFjBZRN2wPiD5j/MCKebJAQiiGeEEIpyoSiDVKjHKIUBuqGgH0qa6YuCTsijoxMShp4VQFYrPSz5DVPD+Docky//dKL4F6EQSfCXvdDTIWu2GVsvbFq23DBDQfASoln2BNXrGuusK0tR2R6WzVB08MwGJ0Rwm08+DHUIDSed+JNKNaWyXsA8VfYNk74tumxJiK9MUkViWPnzCxHM3W47O5xC8y40qsAS3STITuAy0y7xPgUSHiI4JYIf0EMP8wrI/xsvFWmCk0bbcMV9HvroiTsRDl1gF00aXdx1lxWHYfOeNmbRRVeV21I6Hwlh6JXi4Qj2G9M66sA5uMCERwytd2YdhgRPvvjbCymQgIRKPiYM3uyGUwAiGbaEY6BsZWsNIwoOK9KgC3ewQxG2sEXNbHGzGiQhZznjURLWQUIfaSQiRzuI1Io2NaMh7UdCk+GQShiOJEhNJMIYBKD+ZZ6O7Ytj/AKZ/1QhFf5QLDtJFCBO0tQoGpiHMUWEVSpO4jHcBFETOqiYKtL2izioyHBlkcqymiUUSHhIZAGqVFL4JYytcUwKsIMVOlLhIFXI61/60QHHNtY1JLjvF6FZ0XUAof+uO0llbVhLixQYtiLvDLKOeilb2himF+68MUObyATexscwSJzCGc5g3ygj0IxSpqJECevWt6LXylVGcETSEE1oKhgNlumie83an8PqNT50TQuY1BIm+0zJSzpeA2yFjAPLRHSi5hknGqyQxikapssYrAgnrqukLwcoLWDehlqNHBnCHlg/A53sgRF0hxP+oEEN1sxmZliBK1wBQp7hyIQ+exrTVtgjf65DJAoJ6JCkBsMXIqSgHVmBP/s5Tx1AgpTnQZ99UoLAQGazP2MCGxdZBDfQpGlwg8vO5KwDUQPuxoAnnRZH1xPIIvotQDghIxkh8cVB3sRwoNGSfXbT0z//uouQGZVKE0nJPv1oSRNuxI1Ss+g+uK3oUNapIzoQgUerqoJdqeAGu1ixIlWsJzuU/Goq0EELIeimYx5bwCne1dZ3MesHP2hGs+LaLFSOSJXhYqUrXXkcWEojPCuqYAWzJw0B/k5/wOMBD3TB1tAQrxnoMR7mENssAfYKMsgcpC5MlLJnEica0ZRlJ9VIx+uIhmHoQk8wgykFlxlsQBH8rHESRpwxOMEGIQiBOzfYWyf0www6S8IHd8azbriiG5vQ50EZWkJ/3qifCBVoQWmIhKkVbYUVoNJCs3uQFVBjBbTRJWxWK0zWgmaQd1KXdT7KnVm+C5nuBY2vMLtenNgG/5zSotZ9OuneNMZvRegCXn9PQR0D6yIOAKLjfr0pTEhkT403BSn4eJkKBpvPm87wpCDVpeAEB5iX481b8qTJimjgQpYB3vBH6Vi+3mB4WiVmxYxn/APL2rgZp7BxBChYP+Vs68d8FbJy1nAyO6SBgkkWTho+2bsfpOIHOg5NW1MBvFJGdjyiDB7wbgyOSiGTjhWEgzSopy1whVYa25txaG6iLjeLhpqp4MEo0RNZO7s2jcz0sV9ViQ1FZHC3gX5nPG1Yg0x8MGcfHMgHw5GMXvSCHd04IUSw21wd0XMF9DhIPvvJQh/909LPHQQJST0QeriiH9QAlADRBVHySGGysP9GDw+k6WaJvXmWPJgllC0bYvFBckURACaRZG287eAPXb1aZoBUpKIY9HexqDSwgQvWq+KZl1oR4AGSKxiHaoN4l722MLa9iYRmPHkvBrYOgERWTQo7DDTc4KwdomGH6hXSvanlsCowNxHWRuARcKC3vUN7ilP44+ByTjguxixb5KwyyEOWnriIMw04cCMNBBd4NAyOcF3rOrW41AUuulfKHzhsrsHzBy54cIqPP1JdCL5lgSBo5gbU4+awjAa3u+pm066Zxu8yJTEdJtfgvUuwAtKFzaFTnG7MTNC71WA4zOAKRNszhFgfyCCSwQhSkOLRYMiZcyndT1J3BNOkdm7/p5vL9hWKpIRUGjtBNHlcaoC3GXAIja4dJoU7N8MZgGerYG3tZly+S+RrTsWzn+wPKPuOw94Ott8pj2V6Udk772rZIJUu5yqzgpolDlG3C+YdwFOePFg+RfVSXDA3+47L+mN1eYcnSvJ88l2R7/kg39qs2NsVlQMX+GBdRuviI13Ow4ssebT8DTg43+IWx8X0HzH9U+Di+riIBvMgCGSJfz/iDiTzcE62fWoanNbon7E0UFz94MXVxjs+OCto3XIKIjjm1hO4OYejV9pObw3I7P4GqWBY4fCkCRcaRsdODv7OLQJIjveAg+loyw4aABtswAmkzhYEzQbkiWcEohsO/82ers7QVkARHq0XwC4f8iEZzMCflGvT4k5HMsEVqGEQbkTtctC5dJDUqmYFukEGp6QgwoER8kEEzODurE7K+O7kSsnkHNBlNq/wHAnoDHDNwOGTHE/XnizKBtDNIsAZnNCUhi54Ds9lvqPn0oA6UMl62Mr6gm70lC4NwiN4+m48xgMSGO7IEOzbQuMHIC/KtI2a+k6ULA8Mce87WMbNkGyzoIx3fAcSt4Nd7I0SWe87zvB61mXOsox9wpB9psGBpucRTmz6ouERTtEUpcP7wI8Vcc7/hgMUQZE4nO8UrY/lpm/6No7eWg7hoswXqwwXr28AEUzJ7CAUDQTImOMb1udgFGVumdJA+0xM+xLQF3XMGn1xxqxnsDjL/5ojBsxgRqLOFqjuhvzphhZtBNMx62pgBYpwBfPh0bxOEUJgB6dEBjOBGujpg3bQuZSLB3cQ1VYgE3ZED+iOCJOBHXqBEfoh1ebpdwwOyuJqAX3RH55MEZeND58RxShoI7OH/qrM5UCS1qTJevCPruJPIusqe6pn4waQguQwG+EAF7hNeUpmOiqIFeQvrvSHB4xxD+eQ51IB4Qzu/D5vJxmwDk+OrURLe27pGZvyIxmGmnSNrSjI3pzP+Y4sDbjHZUrMehrmDsewlCAhIAAAIfkEBQoA/wAsAAAAAPQBGQFACP8A/wkcSLCgwYMDBRR8dLAeHED/vBmMc28gRIPTBq5p8C8aCoQDAxS8pBGkSY4CFZpcafAYgDgoCy76N3PmQAynWAqUgTAjHIOOdB489K+DwAKEIAnMKPAXwRwC7QidSrVqwRcFWSwRiEelQTn/wAoU+0+ASKto0cZZ849jTIKCQKb596XgBJYM/7FNy1egBax9rVYk2OhfpIMxsx0cTFDaQCAGDxdUeJbg28CYEbpwIRCVQE7/wkSbWkCgm5UACIYyuPpfa4JGExVF+FZFQY6Rav0rVpAxSxYCoR6E8a/0P88FEwiF85FgCZZICobxxNKBg4IeMludm1aqQMAElRv/7NJW4N5/oE2qemNB4BPtQm0u/heHYGqBhQ9+Cyn0vsB6QqnwAib+HWQNfF7AB99+A10gkGwEnTDZQCpYAdVrBCnwj4YEQWjUQB2gkEYav9Awxj/GsMDCCD2ooMIUgexgwQ6BqFBjD4FEEcgZgej0xQggnfbPVgOwBKBAeSmoZEyXKfmPbwcVKdAJTaZVpZNYTpVKk3Dkd9KVJhGn5DJZBobhP5qct5JxVAl3UAKhKMBFIixMMYlAygxUjkCT7ClQNQn+U41AXgz65z97GopQoH4e5IUXU+TARwmV/AOhQfKBBCZPZU7FJEgMVMXEQD2gdZ6aB2V625NoldrpQaa8/zpQfSxBWaZkXoFp0gfaIVfQmSxditYcHDyhTIKNlnPMP4EetEw1AmRTDAB3TgIoJseU4wUmBnmhLLPfesvouAOJW+4/yyY4CQA9cKHNBrFqVwZf4LEknmUD6RqYL1SlIhBHdhzI7XcrYZCkrAVpcMBKZ0nJ1wMD/YQvQbROVXGWEhcmkYJSAXjZFAQJ8JM9B6mzUgMoY5aaBE+MALJAe2qLUMzK9ADEoMqQieidCvX8BgDVAJ3WsgIR/Q+ZZDbb7J18lhWFH2ykF1h7CAu036fwjcoEcP9IzFJcTupLlQ46CITDMGmdIRA0qh23khYG7SV2VbaipapJugx0MEiXEv/BF8kDccjSW1RTtcs/PdQJM6LKQHzQCHz8k0suIEPc6DLl6FwQsjIbpLnmBjmuZ0GDJsit5coqKlAAAhCQL1WcEveGQN54LRACBxkTGNYg4V71fnV/9g9ntKX8L3yb/bMBWipFgSXgmQWvYGWICeV31asKRAtV0tTS4w4D5SmQ6OMj+k8nBgQTyJ4PlNN++wY1WtDAD+Rpv/nyhz86kC8XJD5BjbKcQO6zA3I4BWGhwgzvsiQ9Jx2pPNphA0sWtiGE1eV40MOedryiQZaYQCDkscpdwlKQExhjCrYpCGT+R5AR5OIfL8sfQeD3Dxb+o37lyOEIYmEJQ5gPZkDS3Q3/BYIGNFRBIMEAGcieA8NY5IIKwKCCy8pXPoiJbhJv2EXe/rOSyFmFA2mBh0EW2MEsXYZXJjkgWsZRxoHQAlVtzEwADnS8OGbmhf+AClTUMIUp/sM2aoChScQ3g2TVcApTiAUljLGDUhmiiCMYQTCCgAZgDEESt6iCy/rnw38EIxidRMM/0CCJSwLDAEQc5UAqKQlJ/EMRQ1BEJwsyOZCJrxzV6JEvspEKdPiLFr4Ygx3mJhQM/EMIu3udQdgAxoEkMDBslBVHGngQEPyjRwKpFEHYZkeC7OBwBGEIHLtJTr6Y4DonGYgSBMLEgnCBCzMYgRr2GEg+8KF/A8HnQCYX/4wd9NGVt2gCLC+JSYOEoA8D/YckgOFKgRC0Cf+4xUD6EAKBRrEKrhzCH2whUYO440T/oIJADJCBFIjUk/1TQyQNMQMfBqMKyASQb6gXH5osaSDUhI8oNMgWXTXnH3jA0ghZEsKCqMIgWwFfgZBkFUxATFHemYoEyrjUchaEARNggza4IJAZ/CMWaDAEMCzxjybcIpJ8EGkQBCmQQKJIIAsYCAUKkgeW8CAGPOBBQXSRNzvoIgajWMACeBBXM0BhJUdywj9sEVFJoHIgwZAkWYNg0hEI8R/iqAIFxLEJvaTsGzSdSrwC88CqPFM77WBgyohp1VJQBXwFGSdBsGAS8v/hazQGEZJB7kWeosInAKG1CkkQ4tuqTOAuXDUILYwRCyA1URwQcGhD/zFW9QUCZELsxkFA+g+9HkQXuNAFK/4R3vGWl7zitQMuvIMLquRVCK4Exlr/8dgMyOMfKTCAFMWxDWQKJHi6EUhQQpaWenlKmSBpplWF4haBKGXBINlpGw2sE04ZRDYmKG4ZWYulWdhlINnQnXNHQAVLGGCtQXjsWjOAjCMU4grh0AU4fEGOMfCgve01SI41yIO/YgAHVRhCBvZBX/oGIQhUOPGRDeHCbWQiMNaQLVpS+w8NHCQjUjZITlbiIIFcwItt5HA3XfuPaJrEwm3EZqnuQBDwAEv/IDdQkESqmhkyU2VUOhlvFJ4wA6jMwBLAoG5B5vsPQlMFF+MtyI4JsuNFr8TRA4mAQVJM6ROfOIrBUEMrtBGO14nZKiBIYUEWRmXalOfTCNkDJQYCZoQsbMeoNkmWIWxVJkxKTEoSBTUgSJXZGYQ3TkKbhCWsEzyvhLYCKRWQgGSJYIRUIGQN9EgLIm1BA6PaLGFFe/v6j7zlrb1SQTSOMWPpU1LaEvEcASXmYIZO3U1C1nyFQKwsEAqauo5W0RUMplomYtA6Leg0SKL/8YT3HIQGCaaKwQXiL7aQ7Kh9sXOrnAs6goiaL2KctwY2/o+AI6TVIMFAXC7xAhDEomUD/5lBMFCJyiEYQBInisY7MNKMZghDGPTQQw1g4QpFGISxaWHHNgSCbYMEGpWETrEBls70FFMhspHcRzrKNFSC4NZKCI7jrP/dQQexaSCFEwjXRhsr3wmFzZ7FjMedtBWCxfYfgLvIGEGogXFs/AAbF4UoRHADSAsE1//ockE4YAo5nAEFJk/EsmfwZwMMIQUCgbze/NEMhJFBJ/Qwgzgee5DHMv3zSw9CJFW67mGIQCfILk7gWVIkh2WGjH3ZQ1UANOt7Td1JHMTSBRNtdpPgsSoSFEjwTfIEba7eSRoGSU4PDL3cL4UjDri7D/CugTkQeXJyQIHxDOJFDixiEWwwRf/U2OAHAvAiFyzgA+P/jF/OR3cgIUBIDKbiXVMRJK8Cwb8x/1FXgrAc9C6XAkEQWTNgBZYwB/R2EAejC55wAZWwB5XggBdAHKrAFmvAA/vHdSYhe1aRQUJhbwbha4cTaxBmfG32D2GnExZQBDvwBrCFEEUgK3fzBjS4A3igCj/lZSahWwihEKrzD9PwCDfQBaKwcQqjAfGQXAPRCf/gQ+7ALwJRBlJYBpUwARzAABzAAWzABi0QC61gTzOQC5wHEpLmDP8gaQKBhgUxcwLxDnvzD/HHElvQXQXxA3pTEP4wEHZIh//wAwPXfgGoXyPAeFJnZcTGFvfQAI/QAN+AMtH/cAZPQAmVEIGJ0AKUEEmYKA5+wBcgeG+85iRUllql1k1KiBZfwIMaKBDXwxe+1hcOQB7yFiY7MIuYMCMWwAKTWAmUsAqr8A8w8AJ3UIonSB9wwB2FUS2qgws48A9dEH1HeADzAAr/gAy8QFarJhAvlAt80Aqd0AK8QAm8sA/7gG6TEgx/NgQgYYZkOH94gQ0MUXkgMX92KGlqqBMRsDdxtRLLiF8p8HgpEAyxwAKWsArDcAOLiDKN2IgNsAbkQAS5MAIlsH4RGU/pZgj7wFWnFTEg4QP/wJH/gHc7ZYJwl4ptFFQkaRVssDzDJxSVkkKtWBCxgDhOMjvssQMqQCm5/5gIzLAKXHCR+8ALAuGNF8kMLfAPuxAAjZANgAAIjSAAk+AF1uIFABAAgACFyuEApaABRTh98UAH/xBdEIAMEBCW8jCOuUAJ+9AJ5tgK60dWGfAPhTAQRzAQNmAQ6hiPCOEPb/gPefgP7GgQeXVXd/UP+agTcZgWKVBSJhUMfHB+sSCRkBmREWkMfGAJKbAPQpYBV+AO7oAAbJCRCAYCCCALzngA03cAeNcFA5ALvEAAEuMx5VFadrSS3NQptpEaAOB8J6kZ5BSLH/RBVfGCEfiAk5gLsbANcyAQdQUKJJAHvFiWPcR4oydPalCdU8BHiKQGVhCRwdAJ1SgO4RieRP/GC+RpCZYAjpRACZ2QC4ZgmczwlisRl/B3EGWoHZ9gEiHQbuxQELbgDLYABkYgEIrQDeyoXXyBjm+ZAVmQAQxKZN3JD+KYAdugoBlQCBS6oBnADxSwEQ0wh+HHBt/HAAwwAEqAMg0QDd4gmg7wCno3DHSgDYdgT18IjrmQH2qUGc5lEp0oKyloEi+oJLYBGdjjAlLDEiA3FekBmgKBTiYAnGiRCwt3AegXBRLACwiQB105EKAgjQOBDHApZCCBSpDHeWA6jfzQi734le/3lW3QpQQxlyYhnwLBCPDBEAyBDeT1DweDpwIRA3VJEH/gDPvRXjN3D2OgCIowBuzYlwr/Ig9Z8A8VmgXbkAXyYACdgJYZyg/ikAuE0AO7oJTFQADbsA2zwAmmqlWz8I2UwAeDaAhiSFIpkF9j9ZOuug+UkAsXJxDYxBK5ijC1CRJEMRC72qMs8QbWlBloV0ZSU6Q6UQlHGiwEwQaisHaZUSmC9w8MwAmLQKRR8wrzIBBcKhDI0AaPihCSh47wMZdwShDl+g+P+qhxWa6jQIb/cJcHEQ58ShB4yqdJwhCE6o56OhDvALB2+g8zN3P5GhjrKhRiYBDr2rACwQ8t1rBwSqmRuqAYOgTbYAC54C4LB3belCqc0Ey/VzVbyKxCcaxYEoMDkXwEgYoI0Xt9gQBKShDG/3oQJbubBJGRI/oPLeiCgcAFoJAHXmoQkqcThQCxQrGmBbGwVVGYJgG196cT47ZjbIgZIGUGfwCH7PoP9wUSRWsQXooM41oQbdoGEIC249oGbXAELcYPR3AEGTAEgjMQFvYGF4QwO0VsOlGz2AMeH9tB/nEftqMTbqCyQrGrvTMQwliUEHash1MCLDBVKmABb2AMCLAKhSCnU8G0WRKX/TcQ0VEQUpAWUosQp0tO0dWm/8C6A7GmYxm7JBC7sYsMjEAH8fAKGpac/wAcTKQQ4LQSwqizBoG4cbSKmDEXhYsCKEBhVsE15EQ9MRmTPWC8B+G8/8Bm0MuyLuABbwZUkf9QDOQgENuwChLrtmJpFWJQtFnAuV3rtAXBXRUgEKVrEhAVAfUYAeoYA2ZYmKnrl/U6EGaojnE1v3GFBAuAwPH7D9xlEKybtq1Lu7M7lrNbwRBgwSRAAumgDcawC76Wt3yxCyBcJtSRGS4LH9YUBRYGeMELEkQgFsHKMQdRwv8Qw2iBB7vQwr6HGZEQCY3Qw5JBKiCxiWnBAoVjdgjgAQiAAKHwClfgBNvgAS+2DXF7BF/7D2eqEyQgEGuqtAiRBXErl4eFuoT5D6NrEP5mEH8ZtWfYxmpor3F1uoV5xkLQWQJBBlfgpXm8CsiwChe8CiQAyLy4DcyQWSPwU3LQenz/UbdV4Tp+E8N5qxIenL1CocMvCWE5SLwCobJn4DwGIRJQmGyi/A9qgz0lnA2NkMoXgQfHCgLYhAcIp7gkdBB4wC+y7HYIIQ4gIRIB8AaeIA5DwIsZbMGMkMEXfMwTLJZsS7ZuG7fyUAhUXAgudgWFAMVQXAinx8BmjBmDABI1YBKw8A/hLM7/MAiuQA1XAMbyUMXN3GJnKwZsy7arq6WrgAOBsAsgYAx3YAw9wM/PEAggwMpR4DpYImqSEVwFcUQCocN+oSR+g0aygnAGoTY0XE5bNxC+cAmIAGJeEmAFIcskcaMGQdCZzBKEIBAKbRGNAHEbUxY0cDjAdhAfMFch/+ELHi3LzSGzBFEHBVEfTAlsh3EYjUBHIEEDJLE9teALKEABc6gHwlAQ5+AM5/APSbACAtHNAzEIuyYQ/dAP1DDO4GwQNVADOXcOUw2P8Di/IGHV5UwNZrBOZ5DS4iAOV6AAeQAKdJAHeTAHeXDMYQkBV0ACgY3Mf1zMdAAKq7ANQIYBhEDTAsErJ43RcvQPItHSJhHKmhwYt1xODTYNe2ENckcVJjIQ/rUScwgSJY0WoW0YBnENBXHaOrFOmy0U9XEY2xPE9CEQZWMQJ4DUHv0RSoACYRAONVABerAOVt1pgxDO51wDejDVA6EH/7AOmcDWsEDWetAMFSDVUi0Q8P84wEKhjmY41dDtDBVQAUy92/+QeiaxjJdnErXQwuu0EmHAEvvYF7g9EDxdylRx39gT0x79D/OdFs0x3zZtFWd8EwIB2wPBHRrxFhxx0RNBkuhwEKs9FbqxPbQgIXDFF3NxMfQ6EBz+C+gAcQNBAzSwADoQDm5NEBWwDv+g1gIB3QQB4zIOEqVL3v9A4yyh4zPu4vO7AjpHARx+EMbE1q9dELwR0yeuXB51ECIt2kIx33GBCAG+m0yuEya+EguA2Zgh3aUtEFcXN+Wxl8uR2/DxYNpR4eAA4v/AICvhLwKhCuhAC7RAj/9wAr/wv5qQCXZMEHMhFQ6ON//gLxEACdH/AAdWrVj/8AeIKhDaZaAD8dQGceMCId2W7uKUPuk6Mb82PhAwPhAVsAKDkAQ3XtrRsQD1uxKufRDbMxAinQ3bk+BOUuECEQfogOsHUeRo8WTqjTC0cFQX3i/qERh7uOrNUI9xgxI99YkKMnCOYRL1mBN7WBCZjhDc0G2pkDdpsEX68RN/2NOFLucDkQqJlo//WxBwYAdZxhQNYIdOcJgCAXSKYAZmYNVPttZO0As20A3rsAmfXhCUHupJIAwFLwzrgPBPvelUofACsQ4FfxA1QA0rAI8Kkgr1V+5GlRnkDhJyrhSnoOze3kEVQOsrke1TwY5ujhkZsYhLURUN1mDH//Mpl8E7Eb6QesEqVrMG37B1ORYN3zAN3wAHOeYP/rBlBNGXj6Bt/6C8WzTmAvETG7ERCOE1uOAYccAKKP8P0X4QeXgKP8CoeSMNujAib/fy39ANThAOcchYIRAONmADEY/w/2DwAyHp2vXNA5EENdANZpAPgE8QvTD4TsDWML7wSUAPVk0Nel/3CMHwML4ONaDVNXBzji/57UanvZAPvZAM7OAKK7Dq3aWGdriH+EcQA1f24sVUScIKAzdeieYP0VD2AqELUZXxVcEdi5YGjsEQZo89ibbGBxENOdb1A6ELo4ELp8AK/mBeAsEKeTMaP7HuBBFuqO9gHaSbBcEUlP9tEA6+Bl5CELZi/CsRCRKxMYAwTvzGb3N3D4OuHXVRNzbBGcTz/FlXEOz/Kh9SwwQBEPX+/WswcKAELRIGBjDYcGAagg4lTqRY0eJFJf9YDCxx8N8XABf9SBTwr+RFlClVSlzz71HEikQMQmppJ1JDGDL+KVBp79+plUGFWhyA0k7KggPv/Yt0UyKcoRNfqFAZCWLDS1GXRaX4xdpETgNRNXRx8avDAgbTNjx60mEogwkG8vwHd2KHhgQaJhW6ZulSlG4davkHQyInUwZ5ykUgka/BNSgmUuVqsdRFvo8NMpiow2KZyhOnOeXaMvTAsKdVDwVUUvDegnEwr6Z9Wpn/yrIGcw+cZvDbRbxBc6xM1PBJLBXlGlb7N2lgtUnMm0v/x1w5dYdelD8fqN2CMRZ8Nq4WOFAzRdAKazss1WWgB4cF5afkrJJPCQkAVP0DjDIMLoPquaYhIFYqaKmXUFtkvfVSY/DB0ExrKAA8DAIBwqjssui804aTSAEu3LitO4O8SMk5E2lLscTtBtpKu0nKUeGJXNbriKPVLvxng4pMcMwgDjFUqaA1aDEIiBf+GaAxIZu0CJXdLHqgoVSgciiVimRDqb8m95vQyaDkqkymi7IhzaB9clFhRYfKOeYf7Y4pJ86JJsGETi8weTPPibbDE0445xxIUBL/mXPKQQ2S/w6AWLiABin0/ikDtIHeENK9H81b7QmJduEtKlYGssChBSnaoqGX1gjDQSHbsUiyhsbSTSUgHCkQsgMNhGmipYIcihCJaGlkoK8YAsegBJ200iExxTRIir0iClWi4AY6BDKHMBFvCoNabHEgZbRTjg9KpijnAW/lNPQfZd7sbk54tdMuJQBOstSgAPItZqGTAtglAAECKCaSYrwpphhycOAEAb1U0knSgQyrbAeuMhPSl8pS0REsi1qScL0NyvIhKoZq85JBCX1lsBFdDOJSpWvvAFNTlEYaaSB7rAwEuW/ZHdGgnw0xBJgRyilHma0QBXcri5guh+mhfv4HXZWMjv/OIADcIOAUCXvjkInKOFjtJYtRqq+BXGeOikiDxFkpio3WMoiNf+geaGS1U0rWomiudIihjxlc9p+SM817KL5+Ue8iaf6BQ4k7qOKWXZT4qGjyB5TpuSHlBHijmtuUoVq5AqWWaIZ/DKFCjakdmmKEYIIxVLnNq1sUBFVexrC+lcbBNFqaD585QWhpi9KiKNReYz7hhSqvosGb3zSRWP7JpXosmvgnjIHGMGaHyf9h/Z9bKf95hhkoNj1Rg6aYIhhDijbX/dirECcXigeawhg+DAnGmF28AXb/oMJACmiJf7wvdf8YwQyogIYCSkJ7spOI0oz2AExMYgcoONZAnqf/u39YznIq4Z1KNGCQcUykbBIR24b+wYpnSM+FURmV9f5RCYPMQnqhGoGHBjKChgROhkOU4XluNAE/cOEfPTAIZfT3jxlQJQfuS2D7BlI+zr2uCbdogiQKWIWGAMMhf5AgBStSBSoMwSCFQEYhwAhGQ/yjCsAYgiQc0ocmDCGOFDMGAf9hgPhN7jblKAHrygEAALwhEM/4hab2FhTOMIk2fAEhEScZkQ9QBFb/OMs/UOAGFkalBQO42b0a4qOhmNIhj1SJdJzjODBdyyFGAhN+mscLN7hhBCOYgho2Ur0pBMKP3HLiQGJhjFv8ow8DYcdKkmEQMlBkmX3oQwi6QU2H/0RzIqT4RzP/4QR2kEESQ8iCAcRowH/0MYwp4MU/mnAUh0iokhdp4T8SwxVhBA9blmTQfFTGT67kD5a1cZdKOPWPYjbkdxUpykAaKRQsAlQiSlSS47JhjFwYA4gDESYwxFjAf8gufFOoHg/gKZFuNGQbEsGFHVqaEgD9gwcOqUIKLBKCmYIDA+ckYBAMQgUDyMOjDRHHLVrGn3/0BmcW+UIR6fkgVwnpn4erlkQc8I/LpORGFJkqg0BZmBoOxFkpkeRQ8EChf+xikxJ1CEWLYYxYjIB1KhiaAXw6kDZKAhg2lYQbhWmMYCRTKPB8qS4KG9PVjGIB7tDrP8QYBANsw/8AdrVrEIIQPypsYxTSS95QPqgS7kWkq07K6ivisyu2UsQBKawNRWsDiJQc9B+Yyuo/EJvavJ0BKvwbgRUYaAlLmDMlyDAIK6Z126gg96QrMSkPeLCADjbEAH+EbHXtGowR5GKlQMLtUoM3WpRcwCC5GKGu/rEAiWgobzlYwj+22l34TuSqFSmrSvL1D6YVQRkRPc1VF3oRqjDRIrUAgRv4wLoZIPAfaHBsEGRXBeGqRBczNQiALDwtmQ4EF6y4MHKP6pCWHWW5E+EpdSlrXeyqIRfqZd6DhCCRPJwwJS3xp9miogKZVWQFEvnNSg5wgIq0ZJ7xnQgTc+yQq7ywYaf/wZLa6mkRH06kCP+Y8mlE4aQT0MACKiDvLlHXQAX/UYxuc2yZB2LHoaoEwwMJ8T/aPJCjtKzNI6bIXaULDMriubpoCMQueUEHMyD3QS1sgKD/gbd/APkfMj6tPitTAPFWBrwDIQaRVTJfrkgGD3jwhkQW9GSKyAxsBjES2oZ8EQek+r+qecBrKCJkg1ToShLSwDg0oIED3PrK3HUICMrbEG1wpj4ckIMQVOGLXVQhfj8MBhVSYFODDKEKEUjQOyqihwcJQxh6wHa3/4FtV+BgCHamyGTNbW48Y9cKM4iFNmTxj2Y0CdQVUbT0Ih0UgSQFBxN5N5gKJ7yr7pqID6NF/wDe0FQI3ZOfBenCOERRaw2IQhTxyIMfxIGBDzekI6ABWwscwgZTsGEAnnhBLmo0gxLAjhIOMYAa/4EBKVSAHvT4Ns0H4gRXNMTaM6MADkr8R4mcW+gOVoNc+cAMUQxjrBWJ4UD2cIE9tGI8qJVqk/ZQPZUI0SCyEhIeXE2+B01jWoKoTJIowgGx0W3eQwnrUNzTHpVwYyLAWk0aXlMhgbjCAbc+gA9yLQoGtHMglKCEJH6xPInopANcMAUHQM4GNmhjFpQoQRlmYPkCDgECqmFlRbz5jxikJJ/WdoZB/HER7f1jnAZIQctZ72Av72MVOxHBRBKENjtEoQCUqEQl9v/g+xK8gRxVGEEgqkCmijZkWrTYmFB8ItHnWVr6Q6kyRXZwL2HODBMWeIMFdmABFlDiAr6/oXt70AOJ/cMCX0C4Q34DFQG8EjoG6dsrJH7rduD6Ffv4x8odcoFcaKdWKIESYIISeIIWYAAugDwuiAU+4INW4ANLsClQGAgkmIgIMAhnCD2DCL0MvIhNQC+JCD0O5IEM/MCKoLAfCI1ne7YhoALs4oNZkDhRoIDluYcGwEFTQ5sGUIInoIQW4IUZYIEGKsIGagEd4op6m40ek4jdYBWVWLvpoxf48rh/KAseQYm4Kb89qA1UWgmBsoApUIES6L3eYwZtoKhZWIVVgAb/BZyACegAvAgAQACEOLjDOGiEkOCOibC/Urg1vsuDf7gCCICAbeAFYCC8TviHVgihf2ACXuAFQ0C5GYDACfyHDCgEiyg9iuDAGKCwhgCQ03MJbGiIUfxEEjSIEzSIFRwIFJSIGjAIbHiHc0gpi9isLDCIFkyB//mHfbiBU0CbNRACQhCHWOgBFigB9KFEZVRG9KECXsiAOhqChQkLztChM5iIYRCFXDuAdvixXHOACRgIzwieJmQcDwKT42kSAaiXr5vChrinDbBGi9ioLlwJuxESiiFD3+u9FsgF2eOHVQCFbdiGIRiCSOQFS+iEVkAfg3BA8jIGFZiCagCAAIiE/13AAQVIgDl4BRNINVFYLQQIhAGgA0KEgFUoRJT8B0swhFxoBZhsBUN4tgy4iHz4hzH4hwvEQIrgxJTgpoowgk/4hIkwAqFUCSNwCJ+8iCHIgBRwyk4YAUuQxBloyFiYAaFBoH3IAK4shAzIgkwshJzMhPrigrNBmzSIBBBAAFnYOw3wAVzzAR8YhjlIBHKpAispCFoyEGk4AXgUinrZw7zhjFJRCVXKoX9YkMQozJWokQf5wotgjqayFBmohPEbv6djgR64g1WgAzowCEG0iBQIAhjELl5yH16SK7lCH5gkPEugBIWMTeCawAzgB4H8B2QQg6DQxIpYyn/IQA6cCP8RBMV/sLaXYKVS/IdvsEWHKMVHwIUdS0ow+AfmLE6L2DGJyIIUyMWB4M5/AEuwzIBOmEl+kIdtyIJCQE/0XAUEQAE7yMEG2AIEYAPHWwROYAAOGIAziAQB6E8BiII15IUnaCBD2AdLCIaYjEROoZiNaTshqbV/+CowqaGEoghLaSpZS61jYBMGuYCVw6GpQ4l8dAhMSwnkM4j2awjxYoEoeIFDYADIW4V0mIc8+MzQJIF/aIM2OAJMpAiXc4iaNIgjaIN/2LwilQgcNQjiMgjvlAhNlAeDoAMb4ElX/AffNIh+sIhk2VKDeIede4Tk/IdZtC1seCRDa4jNsoikDNL/i8gCKOXRgdgGrlRIKqCCTqAC1QEq1hsCOYVSrxwIrnRKQX1KrjQEXrBCinDQgQA5iQgrRX2QdQyKCq2NanBMgeOKBSkh1ZBCg8C+qLgnDmBM9viHEq2IJVOU7KuIteAMsWEATuACQuiBzjQIHdVNrmDTf0hSizBSioDSoKiAhrhShwjOfxhFLUUWZNUwl7Ct5ryIDFxKEayIJr2IJdVNW1VSWs3RHG0DMSBSMTiCI8iCcA3XLBgCOvLIRZCBh1EBgRqI5kuJC3nX2ghVsVE4iWA0rtBUGdo34bm+dv2Htaiew5xCBkAABBgAMLKUN/CUN4iCHuADLkgHfvjTgYA2/5TgTYrQVYMASmy1CF9tCDvayYp4xYqgAIqovX9oxYHABkFzgpm5Vq7g1YZQSZVsA2SAAGRoIxF4BZ5tCCWCgfAYCE+xEIlAACj8h3/dnX9wVYCSraG4GYNYq6EomYyjFodQp4YAgaEVJgnlqKGtCC44WIoIzcpgCHlFiYZyiKHtLI9oP/gYCG2oPWSoySFISiadiNmTWYogUtUQ2WhVRaEg1g8k1g5cSsIdiCv9W4kQWYlY0pSgWQgggcidXMmtXGQgAVAYAhAgAJSNC4v4Wouor48ICtb6B9aiu4soinGkjYGlCLNriFjAuoFggVS9iBM9nEOQJTJbCdkdCKmdiP+0PY2b6CQhObKBwIIBWJIBwAHlZV4CwINGAIRriANhqQXP2QF27TO40jw6AAVQIIEb5Qo4dYhRYNy8QUFhdQjFPS8kiNad3ISBSAKXxc2ctVkIaIP7xVnIVcnKHUg6yINQWCnmDZHWPY13/Ac5QImmc1qU0Nrf/UuUSGCDQN2qYAqJ6I3oSYkDNghPkAgaOJwz0RG2/QdZywgnSeBa+IdGGAMwQoYjIKd/KITxHQq+vQhNhFPdhFMMsMCBWABgBdaBeLEhgl8hTolT+YdVIIFCCIRdaGI8WNjuM4Y7kJlj/Ick+drd/VzVyJcMXQmM6WLVkGB++uCJGGEIOQrYyjT/39VihxCmQHjdJjHZNR6IRojef7iEkviCN3iDs6UICh6IDR6KbCAchnCNszreKmgYkyUAcfCEQAiEM3hkFDiDKAiDJjADHLCBLciECqiAZig9ZwBlK/22JKAHM/i8oIAF7LSIWIyKQRgEariCVfhWGQbXIUUGm81lXMZf/OVfX8bZPACFVZA2TyCHtCqJbKwIjEGJznVM1ciKQBaKZTYIvTjV0CiJrJDjiQDjISrilViDvvGGSOi0lfAXd/2HPp4ILJAIE24IfkUJMr6IrGCKbOi0dv5jiUhhh3hgh9hhh9ASihgWiljnhtDnf6ABFFCCG+iGfDKIeKuAGliBnBuI/0H4h1emBox+5Yq+iB2rAXoQhk9uiB9IX4M4h38w6dI7h2aogHVYAViwaFeghi3AmEDAZ4OAD5weCAzwhRQuHIYw6NdNZn4eCEIIrYughpRwCoGuCCwAo6B4W4vYF9pIZ9W4EDc2CNBtHi75pzXojSSjiPUlNYcw5sogu5Q4mTReaoow64GgBame5iAux9OIgwEZiDj4aotAhIL+4AVIaAyoAW2rAD1IAldYgXUw6aFAaSv1ZJVA7JPexJIWBommgEygAV+IZ4qY6H84VbgeCINW5otw64d6qMoAhEFOY4Mga4mQaktL4RTGGCFga7Y6lUwwCL9siGUJnII4R66CYP8hyQa9Vg2I+Oo0wGtdkDtrQARICO4IaLJ/UAV0EAIyYARF+IcpdQhhWIeBAGKH+OF/gN+B0O6GANaG/ofy5grx/jaDyKdwWAc9qIBw+AfSXonaHjCDwOyGyAhvdohBVoksC5ahUGuV0GaHYO2KKJ6ogO6GkOuJIN6gCGuJiADifJaBkAJoOQFImA0a25VJo4iTGYjGMYgJH4h4G4jQy3CSNV8IbwjZ0BKI6JuBaMIz/Qfn/gd0GAhISIUY2A+gEAqIgAqomIbBWYM1OIqvhoMVcILpHIg/YPJ/MIOBMINuSAKDoHIG4W7u3m6DYGnz5vJ/0O4s/4cKEIZuCAcrb2j/CqCA204J88WSG3eIX1CFh/ISLyHZ1Zhvg0iFOMASO5yI4A6NUKlxMEFtrtCSCNjLoFiDzkv0idhw8NIMtvEYx4GKNNCFIle+hkBxh2AFGJ8IlTU945K7YwFoh4CK5dnwZOkNO4CKlpENLJGzNRPpeEPBEteSVk+DZJEQjyFyO7ABKHcIW7AFXzeD2k6pJKiB2qby+v6HTIhodngmg0gGMGAHW5jyisgnYTh2M9ixfErvlcjuJOj2cE8C8U6CJOiGFXj2ZMjSH1jBDHdoh4gAkgaxgeCwQG+ZmZpwHoCEUKla4Yy3d58If6ewQO9xuaNxUl+NFVTZDDyFmUJwihD0/4nghh4XaeWLBgsLCjuvgHlvEiLJ4KA4j76psoL6Eqwg4aSKil55kK2IAw5hFajmNar7B06Rm0wKkJSgC65ABKWyiEBuAN6WKDiGGInwd6itKsGEL0A4ivmIvs3+BwoAFoKeiPYyiFXDbUkHuAR+VAzROkAQcPO6iOqzYIPoJHKeiHmuiA6nDU44WsORiFG7iMIhjK17kEuwgCirjaGeiEXgkY10CGBcCRaoeoc4iRA3iDDo4AkWFZQoVeFR61Ojv4FYFvWQmC+8VJppiRlPx4bogbgvu7yRJ4NohKZQe4dwlzSep8UxiDw2iZPHayIqkDcBod3guiaZArqviFCw/f+BKI6qWo8Oz4G8/wedUA99pYjnSRan74k6iIqrcvzm8feUwGCKyELTr7CL6A1VwIMa+nwhSdsBEFX+Zv0tCQqAGYhXmohO/4ccqzJXcwtrWP/TmJL0K4wHUa9Gm/nywyENBoh/Av+FGqjgX4KBCgUmUnhIYYMGcBr8W0NDoYoR/7Jl+/flH4B/AiKlgbPwJMqBObSkbDlQykCKAte4rGnzZk2KMnEOrJeyDMo1OnkOjET05COBGI4OpMT0Kc5j/zAtNHlv4FWTAf5trdn15NWWEngajalQKtSjeHBySjuwIdx/BWxa4Unkn4yHCws8iRLlDchqAEKWW1jOS7lj1Sb/VRu4uDHKJ7y4MAvkFufOhSUuc/43NHNnPgtB87Q2sAhOJC3bLmJg80Ln2C7jNKCJE9DJrwJk8wzJO2UthbsrHrX9+18OhQdPLlc45Z8XyAqrPf63+N+kgdmtc5fOtJwagaIFPlEIg+hO0gM3C2Rx/OSrlEN5l3fPdFrLFzyTXk060NR7AfI2nFtn/OMGU1/94xM6AjqIUwcO4ZRcSgowcMgU0lUHHUqMecGhbMoo9OFJk6ggAyWHVPKEXp2xV8Jm9rnlG1PqPUiUNSCcNAFmT411I5AooWOcg3e0RGSQTxWkkBI2xgabQly40RhiJ30o1XbYNVaYQBseR6JAhZWz/4xAIlazQy7/QHPTTmFpNhBQSaLkpJwnUYSkTc3d2EVsLgy0yE0PODLQNTfRqMpN3wBZTJ086UmUjEz9qA0XKjwA5ogcYjqQF5gI8Gk1imUpEFopcfnPYZxySaIyYG76YTWFLYbJB2wIBKCfLdkYZ6N2enYcEwLRktY3tXzElD2/vpfrQhr844BLCj7FkkK44Xlsrwp9cFKy/zRSlLRMKYGSf//UUgQQA6VrU0JJ8sHCA6eealOqjh2Dyb2TYAKAYCLW9CpTD5xEYxRctFVTuS5ttpZAij5o23y8BWuWsjyhkFJbHuiqbBjZtjTASagcdexEv+H53rDHsVKxTXi2e/9jSCO8K/BAh43Jqaao/kPJCKN2ecxhswqkr75EIQa0F8oADfQyh7WKc5aTcLnbbipwoTFv4ToYcWfBlncTtALpUNOPCjE7Gsu8nU3WQht0BrFnJ3t8Ek2AfFvUP3FQPPfGOPmBEqID9cCCmP7q/E+8JBY2wgi5dDLFh2TW3PRCTyO2qU2YCiZYlwJ9KoAvASjYSDZxAAJIHHrDoYsnCAB6ik888TrQRwmnNIAxAgGWFtd8n1Q2VHTyZCtnl2gt0JI4rdUgUdzcJDdRB7uGXtotRVin8Ar93ZIF/0zx3D+G6wz+4cEAQwnk/5CJGJlkzmuqqziJeZThh2EyCY0WyOH/q3pfz66Qw1LCBd5kbyER+IebenWwJA2AeH7Shu8EYprjGKeAsolI9W5ylxu1qSU8asFJTIIHY4xgCu8TCM0QpxAqACMYO5AXSk6IKsnB8DvlmN9RqiQQAFiAEHtTDxM2A5T/oQQBvylX9qb3DwIcMII1wdMGoUK8f6BibXy7io3OM5Bo1IRAAQog3gRiwbl1kHo0IKGICpPCkwhsBwIxhEYUEi+eCCAAu4gVChUyv1Ot8R8jyF0J9SiiKYQnTCos0UAAEIhfjDEtSjzKUnzlxOMk8DfxcUkUkpSekyBoICapCW4ehC2BSKuRk2TP9Xg0kFQ0QBfkKCH5BCY+Pf4j/00DoVkawzcQZZzwhojj5RQeMAU+xGJ8hlQDlwQ2glYEY2cj4JK/yjGFERiCCjE8pHZA8oZa2GFBe1PIE9ijkmyZEiW6ONAk/5GwE2zrN2FLSQ80WU6m6ChAASiL7/iEEKbwgRItyEUUUDC2gZxiGjowxvcUQi1dytGPKOnjQqYJx3IIM15TmEEscmGJZ4bJjXzIRQkFNoVgGMIQA6HCc0YKx2mKxhDAEAcwclemh4ZpEjvYxTljlzZcKGRiROHAP4Aam3mexBPpzKBArnccH/iOqO95WU284Y27+cSpnOmCCRSiz5uwJ44CGQEL+JC7HpQwPIV0zj/SJSJ/lQCHNf8rjArSVQ6NGGIGgZDmCNCABhZKIhiBaOMIgkGFkv5jF9kIRDCC8I8q/MMAQxjCP4KBhoFI9h9UqIIBmnCLJvxjpdj8xwxiiR0LoAAcaNtJN9PpJA4I9R+PjI2zAtQ7othyZx5bGUrItwYsuuV4btkqSiQggXUJBBAysSpvsooTcbagISr4hxrOCj41kM97ClFrWv/BghI8Z60mHEEsqhCM8ZpUIVWoAmQZAQZFNCEYEhUIY09yXgP8QxK3kIQk/jHZhQAjBYWA7D9s0YQhiHem48lFLHk5gkCE5A2f291RIeIS1yyiNdvgSSX4NtsIc4ZIOk2SDDgsIOHxaAIT2Af/SNVAoYFoxKsCqa5CcsCH5xRmB+G9xX2BsVgWouS+j12INfVLBWsagAyc/UcI+tAE/MbXsikYQiE+gWSFhGDJzRxPCv6hWENYhlqEjIUJyxGIwJIjFShZMU8YAKCT1DMtvBVx8DAokxDDmShlowXcYmOSoXDxPXQuG37qTJQB/mOAsShreJITSO0W0yUYqIIkqnCLf1zhCmAgg0Js8Y8+nATHm/20QiYtkBAIpA+SeOypyZDfk5A6BGOIgR1i8A9x/AMYGViIIZr5nBmMV6OLFUcThvSPAELPJkCdYmttwlRJftMte7hJO7ZWMeQ66J0tea52ByIBqvwjZf/o1lO4/402OTEq0AKic7cfxIUP8kIghSRfM0FLhU7EO6EDscwo/tGNf9gACk/Z90D2PYpN/CMGPPiHHRYw6ikrBBQCyQMdBhIOgbDjCmQQ9Uksc9J/8GIbQwDHGsD4K5oUu1dvrgkHOibozyDViZdMSeBOUoRd/EZygl4IaupEE+EpkQuzYIY4yDCAFACDvgMkR2QF+w9L/CN3Z1UILlLbEmS4hKc8sAMr7BD1geCCB7hgBU95+smbELzg/1ACrRWi9CBYMwVVyIViBRLkg9uG5Bqe9s2fQm0nAu80CqkkTxqgCnF3qidbvAxUURLFDz8oOO9R5UJesIaONBq6/8A0GSC76v+BPOe5PdC4QGSdknMqROoDIT0uUI96rGtd6kKgQDgkgemF6CK1rIDErK0Zdy1TIQMZSAF9U8CPf4wBgy3Bp1t8+A/QBy9by5Zts1OShm/5lm/nmd0os4dbJ4m7Hrbp80nQjZJSBMgboawzj5Q4UGMcmrJBMEAbGEEGRRggv/3dxkYJyfynqF4gqff/6mUdT2WdQoheSozBArjDEAxZrVkWMGyDAbBdEASBIahBxwnBuClEJLiRFgyKbKyC3vGEEcEZAUjYhqWE6ATIXCiELDyLEz0dVKCZVg2I5yxE9wiE3kRQsg0EIH2VIbzf+w3EESADgEmCIkjCMzyDQCihrIn/ngH+A26VXtQJIOttnemlxS/EwC+IA0wNhDzUHxACw/tZQgVSwjbkG1OwBAAEQDGUHE5E2z9E2/MN1XHsXfQJGvlVhXaNB0/wCKHZRDyhBOPZhBspRB4KyCjlHU0YAx/E0QhQQRBGIJAZgI6NWgyAQwyY2crw1ELg1tcNRBR6YihC3cEpxCgqxMHV3ijMXmPt3gRGICwGARqoQS5cWAbyjcicVssdxbM9Wy5UnksIwx1ugNvkHVHIQh6Owz8cohMNYks4XktYW4CICHFFmCCYBCOOQHjMgCXwAiWixO6lRRRyIhT6nycKRBSeRCjqAtixwjlZ3UnE3QQC4StSQTCo/wEfbMMKHNcuKsQsBcjY/coJMkUv1lKN4ERsGaNCZssfusU/coYoPNE/AONCmAJrCYQnnFMU8MEMbGM3atnu0ZdLbF5KtOMn/sNJpmQ6DkQEYGAnoiNK0l5K0Fcs1iQc0WIoTJwY9eMSMMWaIZxC5IFCHMA/zCH/9CNPQMk/VEIsYJtN8Ja5tQRREqVR6uJC9oo4QVhaABdPmFlKCAz+KMRH5JxsKGOAeGUxaQQ38kIuzIBAAAMakFRLVKJl1cQ7ouPXfR076mVMvqM7wuRCkCPpuURNAmEEtpA2UgII8qMbQoUONAD4IURCnoQHGMlV7JxAdoYtZdg/8GFLZMJAov8EUQpEO4zmQmDmVS6EUT1IPAWLODlIQ+IEjKXmhQWOZbhl45jUCDDdQtCXKz4FJxKgQHTTOREnUA6nbBimcgYB41gBJcyBOj1Ia0kDCujHScChS7BcbOSCUqYmnGXSP/RdGvSOUMXmQpzAQnyNGDWmTTAjU8iggETkP8TWZLrF9JxALViABbjBu7DYeIgkfmGAJiDBJiABElTAJmxCEozCCmBAONwAGUSoOEhCITBcktClYmVoYcZiK6jBCFjBPqQDNSikdv4GRdqEHV6lWbbEBain+NFADp4EgOxgSoDnKt0hT4RNC7rFLggAjXAGEQmEKByABhRpQo7LTWTYap7/hA7swguAQEa5B+PMQCcE30BIgjtgwzeQ4z/4gx7oAT0MhB78w5jWgBnYQE1o2k3YABlAKJoOBGSJ5FsOREjCogHcKZ7C0ZQygyxgjYAwwGtdRmimRaTERrSZpneehHsuhE8NhFOmBIDM6FPEnMhBhXw+j/LYRFUhUCjdIGD+QxcYqQa0gwYcgChoQCjogNy85rP9w08KBCfIgRLggQVEQVt+FTUtBPD9AwUI4zu8QwX8Q5gqxJgqhDC6hROgxLAK6z8Mwg2IJF0qBE3iKbVG4Axoo8ysQgs2Q6J263FU31FppUIAylO4RySYRDEIAM0dxxT1Sg546hb8gwh0QSk4/4ADdAFWvUIo4IAQ0EQlFarZ/AMbmAIbDIAnQCkviEYJjMAMzECWCcSuCgQFOMMpFCtU/EFawAJKwIIZ0BpNosS0VisltkJzzgAvhCpOdEyGZdgeBAvDVCpG1uF7ZJj4HQmODmUcKkR93myjDMZNXOpJdOdJfAGEkesiLNBrCMRmiFsiemtQCIQDiIIokCqRHsArbEMu5II4IB3gKe1AANUibAAbcAIHFGwUxIIfcGTDzkCaPKxIPmw4rMA/9ANKNNE74EQfcBpUHJwmoETRCcSdAm5jiWwE3uOHGgII7ixK4IJRVcIFOO4efA2idC308QZstKpAKG5K1IPcooTiyv/hSVzMYD4FEMBntkFFVLaEjTLFRf5JoUHFFxQiUyhX8/1GGpzEWuCHK0RtqfqAqQ4DNLRbLVFCFRxQsc0Ca43twLIBA6BYLDQseOXCwx6BMf6AP/jDPzTRSUBAA1Yr8KVAENzjtfLCKiQeUghENHhCAVRCLlTCHjjueaQCHIyCEvxCk6UETVzM/vDNCg5E/woIdtpggEDUUWjvQBRjS2RYmlSCfewfxpwEJgCG7C6E+O0ACDzqQIDQTeTiSZDrQoBDMdRC7cnFUv4D5qaEFqVEjB7OP0wDfjjAMBipD2hAPHABb3bCP7QCF6LnQCwBr1TCBHAAAyxC2bKBNiRsCbT/QsO2QgpQXehlrzNkrxT/AEvWxN3+qk2QAk+sA/r6BxfzRCGcmgEA352iwZ6mg7NAy1CERQN8Q0RMwxmsbyWwr+NSwi96aOPcBeTxyPbQoUBQrqHWBKMwheYKiDJ8gXrWyf/eRLsuxATL3A68AQi02YPswJlIsiT3AHc6Lk500knEKKaswTSYQRdILZHOcDzYYlOs8q0yQRmUQQlcwAQwgMGUbcLOAEe2Qic08T/kG3oasDNEQBQLhPYekAH/w90qBLe+h6JwURKoRpeexMH5Qykig2ONcQqIw9pawhxogHzih1C4cUSIczTEcR23QAtA7wxYAcPyQgvMgkBAHvpC/1vfpGhNRFsAo0QszEIjHwc8o4QX2QQCOxFZpoVT/MMbRLJArK6A7AAmRPIO7IAFsID7zjElPEElyEDfpYTDGMckfMh23O7DOUApiOoBdMEqfCEOC8RBD0S78UEJzMAT+AEXUAYStwIfBEMn7EMWnKcU/8MwV/ETU/FJ4ILtBCskPOFAHFwxt8TBKbVAJAXA4cSTpQDwwdEMtIIIiIIsUIBQRMQ91EYbR0QDkIMfpPPaLsG1rvUITAYHxKYfqJxNEGU7AG1LpK7THkVA80Y1AokH20ofn4RX1dY/uJG4tkQKt8QreDBK3MHuJPQOqEAJOO4cU8o/aAMEcYEQN2RD5P/N+XmLlowKkZTyqZbqMMQDCCIDP6SAJdRWK5TXDGxGK/DCPigxLs8AGliC76ly3bZEDETxAQWrQmCD/0XnPwij9jbhQjD1T/PEOzwCl9rEw1o10QVDYPFCOtzAOzRAWN/DPazBCbzdoS3s2qozwz5iBnBBYAfqSUzmAfiuDzjABFSCG/CwWVjQCThjSxRyXuNEQQeJC5hCgAOK8CbpP6gAJtuEeUKFe1BFREf2ZL9vJbSANjADbQ9EBjDDKmjDNviBH7jBF0QCLaSO6RiFF5DIdsRBcCTAK+QBSRcpkdKwUArEKkAAMmQAMOSCU1yAaPACL6xtTGfUPghETytEsir/hMK5xG9DtUsEdUpoL1H/AioWXCkScyYM90LI2jGfBHUbgEmVQC5UwTMQQCyQUHk3bEyn+drmAm0LnzjcAhcwr0LIs+eAAA4MQwyXamnCtwMMQEOcQUCCBkz0N1PsdWx4KpAACBu4ACdwAgN09km4USv8g9DKBp9wZU0k9IFHuEWTLzPMgs+JQwb4uI/rOB/wQSskQi4Ywy6EjgB4yImvISBcAg4oQAIkQBdEbUmLwjBsgwesQo1DgLAjg42r9iqgGKqfOm63G4D9QwZU6HH4Aydi70kQNUr8ARlIGRgIBCn0wkBIGUoYQVo8GYangO+lwHh1I8PGNrs3rDFk9U77/57vDUEGZMEN8IA7xPlCcMH+RkQaBAAK4IAolLQG4EOpHvwrcME+8AIhpAHjAXIIPUg/J8mPxsa6YLCACPiiv2pNVHpnKBc8QMVkP24lUMIeJMI+AHvE/QOwb8PCWwIldEJ5e2h0EZIfsW0sEAIhGAyw3/orvEI8OMAriIMxBAIXrAIoADsE8AMvWEInxHwnvLYhyOk/NPs/QPtAOPFJAPdNJANnfAK4L0TY/4MWa/E/jD1PxMC2wymc/t6o4/Q+WEIwUIJV74O8Z0G9530hZIATuANNZAICIBsCMIAfNElE6EIkvAEXyIKue/MwsLwl4HQrWILyPUUUmYtCnKhbcP+CFaUFohtKnRUBJXewq2Z6YbdEX3dG8pyE8EJGIYbY48Z+AcBAD2xDPPxDxK38P+RBjfMDP2SAl1t3CZUVIdV8dEXXlGZ1K1ACJfBC8zd/Nz6/81uCJaSAPPBDFtjirS2EPCwE3qe92TFFkh/nQPjHN0y1QrwDNnSuQIDBGFR5Wmz/9v8D3uP9PhjCbDNDFuD9NgBEhixZ5A0cwq8KnAb31mxBwGYRGw6cGDDwo6RBmjToAoBA8OpVulVc+MyY0YoPSkq8/u349xJmTJkzadacecBmTp07ecLEBBPPFwA9dar4V+Sl0ZwMJuSs9s/Cvy81Z/1bBPNqzimBZPy7UID/6Es2Mp/ENPGvS1iYU2NegHkhF4seKsTRmReThM0UMQ0AAxbEkiE0wYKNKDzDcKtOnSw1tpQixbZtEGIia9PmnxhkanlGyOls5qN/70b/Ey36H65/2GD6c6ao5iNsjx5t+gcbzD/QMUnvtMEzg7wMhTJkoGIpA78j27Jsk4dMXBULgBo0gONQIqeJDBb5CTRphwpCuQyNMB8sCOR9uYKd5LOPJcyoL13Or8mBc36a0IgGqulfvwBhAiKppf5pyqZlwroqq51iCZATAQOM4gUiOOEklHnoqAmCI17KQKa9XhqCr5jk8XAztTArxKYsZHLxnzFk2g0mz3JiTTXUZNLx/x1/HvEnhnVeCiGEGFhL7UhcfGTNH9Z0lPClgf4ZiKCYsjgigxQoIS+XXCzhZQhexOGFCy4k2wZM8vgwxEtL/kmBxCyHgBOyFPYJjJdEZvhHKc4OCdCHlzTQb1CbcrFvJkShpKmURR3VD6yXCuBjUQfUcqmnHvw7hAFOTHGBEwXmieefPECBKcWZSHw0Jsww0wlGmOR5iZEmarLxUR1R84c0XFjDxteaesvPlfxcPMJDD18S4x9+/kFGDH40E4NZZo+YdUqBPsxgiCyL4xaYTnjJhVX6yo0pwnPPnUNdAa/iJCsOEskJQJgKKAupnK7Cz6ZGHUirpqnylWkonvg1Rf87TrZRYMO8XrLsH+JAfEnEEGMaIotCUqWsJ8w8ZPGfiaeMUtawcI3hnxgiCKHc01Iz7eWXjozJGZRr+k2mZF7ML9VXX8KMn80ws5agorP4NgUqMjj1nyfKMgpTnhqUj6hAYUpAJ+44GKsnBf4BIaaodUq3XZ4YiGkAR/Eje6cLvvoHrEDeAPuFsmHqgNyCBeiJXJgY4KAiLtx4441AtqEDlCuejTg/kXnieNmZCorVxVhrWiAmXF/S3CYeSoPpyHdm3hFmmT+HqRueaISJkZlcxFZZZmESQ9lUbWoDAtxd/eeINo6g/QgqM+BlGxNeSeBsmFTY4Q1z+ZZJUSgRTP7/H35rEsVSm8S2O8Czp4YSAZ2ajwmGl9xyK6a6BRSFe5oQbJ5wwsWZI4+d1VIW8pkoIwFyZPVDIiaYk8nJaiKCmIyDJv5on1qwxSzb1cRnNskdBChoGWQg4wgY5Fb9unAWrJWAJl8AG08mUJb8sC8s1KvIAm1SPhbSZCgF+wcgdsIFmNjQJuMjiwz8E5V6ySR8L8HhTBCIwhf+I20xmcouesACFoygB7lgxirEECeS5Sd/dgPgAHUTFp29xGY8YQQ7jvgwzlAmfxRUIwV1BwFk5IFUnNlFTwiRHwS+BGA6CeI/qKcfHZYRkDm5Q010aELlvQQFOkFQTRpFlABwr3lO/4TiSwrmgSuIAAKrKATIAjkTZSnuH0L4B+YEKAWYhFEnLNvcKP/BuQAJsIxolCX/KMg/W1YQFHRYxT+yVxMJyGRve3vJLhLZyXLB7x+7+GMZ5aCuNMAhJjR8CQEC5AYZuMGYMQnAI2nCgp18wCaDtEkoOOGCmFwhFNu4wiYxJpAryS6N+vPkA630EmzJBAlb/EcFWFkjokTAGTbyDI1AE4EY1CxlKTNoK7n4EimQEiawrIltaOKs3f3sJWusJQRueUs3gmIVBJjjP6rwklf8A2sggUkSc5hNl8bkhzApSyy6Is5OxgEmqpnJSNWCTQH9aYHe3IkfvtZCcRYBDx9wgf8HPMAJDyDgqU8lAB4i0QhAAKIRkQjAG4yRiyFwIWj/WAUoyFpWUOSFBA7LIkwsd0XZDUlGM1nAQ3eSG1TOBKFhKWgA+wmTTSxAn/9AwiYoOjuhIWOCuGPjGmnJUcem1VR52IYcxLnMsFiWJ3WsSQ/UUsyX2mSEMPHpP6Lw2UXhgbQP+odQQbBEmfTtpZ79RzPVMkihEmIbCNAtAnCAgwH4tgoCqCpWixEAX3DVGOIYwhVWgbg8rBUvMXnrP+5JExdxslzh+AfOZuIZV9LElDtZQGFjZBtN0GozF7ygG9mLWNwhYxUQICsJtoEDcchBDkSNiRyMoRMD0mQuNOGmTb7/wNNlNq+0YdkFT017LiLABKisguZMAGRT1ArAFzG5BE9o0GCYxNRuOLhBFZ6BgCtshjj/sOI/IjgTh+3EfzuxnG0AGFhWQnRR1HjJCniiTyGJ8iXknck8SDAESQBDHB8gcRQC0WSYcPYlUQABavPz33Lpl5oxmeOGYxIpDy/Kpqy6gYAmnBNPnAEmGTYzlLMZiX804h/HhV4y/0FlnWTYzv/o705wEJNiXOMf6ABENrIxhio4gbnIyiB8/8G/nDi6gm2YLnZhFDzahSwPInCHTmxsk9XlpwYvGcRLXIHof1iZJ3nZzCrGOoRnLFgAc+tBD4zRA0/Y+gVTtsmDNSwT/6+9JBRlu8QuuEzndkUYkHNMsEzYci5BSEi2aOYMiHmiPqKAEyaebQScY0Ll6NEkyzx5BpS4GcxkBoIAOGA1HfLwCjo4FxSRTesqSHAFN554nYUggw0oEI4tZIKwFajAOSqwCSe8RKLqCrVORv0PWDicGpbchqJ797veiUHSbbBgYtVob8TGexsECESta/2MQIRWJxjGMINjEux2EdvBMKGtZiVEgzrohOXZTENOqgOTBvS6zsV+iZs5s2E1xyTcNtmjTShAE2twOwB7G7ZMagGTps8EC3Gm8tH/geYXLJvpz4ZJHHQxw6G/ZMDegIlmNXv1l1zCF5e4hBJukAk9VP/g7i/h5+oqUIMVDGIQ2vWrTMxAxpo8/OE0WXji10EPxycBJjVAPE0AT406oOAZZmI1CS646AtqnOOIFf1Ga3kFEqwisiEnBzme4XarYwDcNfGATQJA9H+onSjC/HKcd68WTUgjJ/f4x8+H34A1zKQY/6i6KnbOPXL8QwmO4nZMqi4TVXT4H1nP+j8wQPOqJ/8fNJDtP8ZfE2nCZOdZfYn6X3L+mGAAC1iIfoZroeZdhMEV3eDnS3ZzjpfQg8dmAvD+wRX6gQBnYvL+IQAV0OFqIAkErhnO4QecoRn+oQJpAjT0YB0WLyYGgRqKhfxK6h9o7h8O7uD+gROugLnqawj/zqQFt8EJcGAbhsC+xAELEgwFaADuZoIQXK/64kwEdQJsUIDBiG76PMwTjGnDyi+bju/nhO8lpAEQrKEnaIgKFyUMZCL69CMbwuIaaEEnLgH8YkLaoMT9ZIKGiknsdEIJAkEJwuAGtkAY/kEPpEAPUgcmGs4DB6EG9EAY6AEWEo8mYKEG6EEPmmE3EFEt/M//KPAcmqECnOER/5AA1/Alti8myOAf+iwmSBAmki/5RmoLge4fshAT/+HmbIITiaIRiuEIYSIJ1eIUjYnrWAVsQGAUAckJ/wEKreMfcIoncMr9FoAJY0IVXiIMLBEVY0IH8uME/iH5sgEQwDAmquof/yKBCoFvJ6jRJpoRSqjwCttPJoBMJrhxCZUABQSBAmqgAoRBAzWwAlYgHFaAn8JL72RC4AYOJvxvH2cEJj4NNPzPHimQn/iR//qOGjBACbAPJlJRJ2Zx2v7h+WpiDGuRKMaQhs5QJspwDHvvJcCwForBIqEtQMiRM8rsCYfvJcqsJ+IA0JTvGY/ovJQRDGnhDDMyLHKxGKpO6BYFGGOi+V6CG17iJ1/iGGECDGmgw2hACVZgBRqPAO3O//avJviJKvePKmnEIGPiAjHwHy2QJvpuBTLBKRmSJlzvAP/BHWJyJ8zyJTrMIR1S+f6hCwMkka7wqjRSJpqxLj2yJrgRSv9kpBj1IxO2ACbYcid+jvgCJBXesoy8sWwQgS5hQhUQQTIlZOeCUibgYOca8yUQMybQ4SP/4RcoQAScwAnMIBzo4R+EBCvxESZcszX3CSaoUi0Csot4ogKSIBwekB5cQRB+0JhESQhMMhtogRY2bYFE0y9hoi/VAhJsAjQfZQ7/oTpjgiWP7/heQjH/oR7yozMXRQqO8Sgf5aqKUjPDQjRpIQIu87tk4rxkIjPhwA5YcibKzjNX6R90AQ5Yhox+Q7sWLshmQkju8SWEpEAroEBhYg6tsjZ1wjYhdDed8v1gwiR34hkB0yipsRZ/4TJrwhs1lCh+IfxeogvRAadckib/Eo4nBBQmPlQmntNRsgEdylNG88MtTVRAAssedWIaYGIXuRNKVCE686M81eUnf1Q7e4I5M2cn4nMmngmaouEfWMEmWAEOpGHnuIEV7GAFnEARbAEm/uAfzGABXwIPrzM2aTMmFpRNadM259BNGfRNa8JN21EYwkFAAcjfZIJFaUJzXjImSPQZvesfjtRuyhMQRDMV4uA9i1QnBCEToBRKyw5Rm5M5TwBGdZEmurNcyo5LtTEs8vNyZqJIL5UorPQfTuEHaoJUSfVPc2LCtvMfaDUaoAkOchUO1sDgFCEEyPQfxPQ2/sAMnIAazlQmWBPy5tRAY0IY3FRN19QmFHQn/9YhCQaBHqPVFaTgBKYzQJiTRGUC0CDBUN+zXJqUJlKBVG2i0xZIFVIBVY2JSqtUp2qiVXWC+GjVU/ODVmNiXmHCDl7iX//hB04BJjwHJhozOkEjvBQxYQv2BzwHp4ayKANWVWXiG35uDepTG6Oh7P4BHH4RJnQhFVihZFUVV1wJUkUWSGmCVtcgCZwAWGPiD2zhN8wATf8hE/4B8lAnCWogHJKhF0ihF5LBDFKnZ3NCSIQhCazVWedQyGriOpP2WZuWTpMgCbpBx/TASofyM3KTJnAqZP+hZBvTMz+WJlTGUS627IryJXggPz/WbW2iR3XiXgVkXX/RM+dWP1dSNf8ClifyViam4RvW4BteYg2ehCj61Sb2dTFj4nF7bjuN7x+g6RFYMmAViBWsVDVw4RRU9RSolFV54AcgFRJ+QIFyQhdYYWCnYVeFtFZb9iUC1g6kwUpZIUVZQVSBLxpOYWXvNgI8h0tfovmg6WXztQEWAAx8NSZsIQTCwQy4q2d3diYgLxMWrhvMoHWI9iXyoRfA4A+6YRPWYXyt8x8oKglY81jpIWllgnxfQk0hD2vbV01XgLt6IR9EgBqSIHVlolU94277V25jQhdWNzWkARcA9x8Q9iVa9W7tdnN+4ALZliZ2ThsZeOzKBlJZ1WAb8167kiYUeHhlQhcMtmDJdoH/yRaDTSMaWAFtqxSGTcv21CIO8vUVO/WQmu0aa0L3cI8yeWJfj2FRHuAlBIBvZ8KcYGJeH5csZALbeMIPNmAneE0mOkAm+hUMc4AniI6JuefXAoRAgsmIbUK/mnMmurOLew0y/yEAhDgsXOFJ6rV9jKhddM8maHWGiUIvX3gm4kAvXyIcfYknJsFRvOAf7HgmriKJoUQHlABV94ZAXkKK/8FrvrgmrNiK5yUmflQmtGBAeiKNy+ZiiQKEQEgm3PbBytiMo8nnYjcniIAE3cwCtEACyqcFYqKRrlgljWlgWEWGWLYmbph49WMwZ4KGuO2Is438juiXy4WW/6FuNgwR/0TVJjpgki0ZFSxZJuaFm//hGdegAX60AX5Qi//hEhh3wGCXJzz5iH4pJvpEJ1jqJazNL8F5l3fCIY8Pka04LOSYJ9hMLazmJVAukIT5H9KzJ3RBh//BjWvikdKZO6XBzSD6iBo6JrZgEa7CFP5hkWUilHNCOGnCk9kmJrT5JTD5H/i5JqoukmOiX9P5o3lCQXSCXWCCXQxWdgf3JdyZ52LiGnx4lWOCChlXQFwILXgJh9VCNFGuEjyymW3CzfIYoQXkqYv4kHk4qF+CbIhaJwxpJ4xikU36H6j4bmBCk1t5Oz3ZCl4CD9YADuBshu2zJ8q5hWCio9ViXpfAJqp6v/9mayccoJd0LqZnQgc4mXGBQK9zAh5mImD7KF2LCp5ZaOmiNJh1Io9ZaCoEIAA2LI+5oY2zyaJpYqNhYvZ6qmleQrUQFyYCABNa+q5jwpy8LKVn24qp+Oe+k6tRS67z4yf+ga5lIrFjAhUCJEfLJrCzWkjTmKd7GmD/YbJnImQJuozkGTsB4bJrdbCJgpCvtCaOga/PxZBnIriJwhHCorRdapJp4qxDaSc8matbmSgi+yVAaAmMWids5KOnobg9krp7ogzUgrZ4opd34r2JAn1eqL+Jt9xWuxHsGaofZY0LBAAoeoFMuVy+hyeAWlKoDv06UhleAtlmgj9AuVZ3VRf/UKCJYoEFSoAFoiCRAoGzomAEyI8GaIH5pjomsu7D1eK1kVsthgiJuIesYUL3Bpx79uAfqqJ9GCSpa+K9rTssvnsnFprI2TiQoWS7/wGEjHq5oWS4YyILIbcmDjypuam3/2G9w+IQVNoTiAkFAsECVAAIgKAaniImslyGqgEAMGEHEIUlmOElFEAbdjirE/xRsnusvTVAqBsDTiGNW1onInxgfVw/fu6P4Vub8sPIlUgnpLwnhKpdXG6B0nwm+qgsuDkXSmAElKEaJmEoCPnVGRomDFmIFURBnsLO/yG8Zx0mhMoo1OAfupx87FstPhrUKX0nLPylju+5kX0mrlsc/3uaiRHZX9WCymWCwhsMFUQd072zXJpaJlChpp2b17ApF0ZgCnadJhqa3cPCC8phEtT9JSYhKsqCBX7b2YU8J/77Jbpi/QrcZWeipemZJ+oBNYA836M0SGHi0gG+bBB9gYQYADTcpdbapq/mi/9EBlSgHI7h3WEi13M9J2idJ7zAkLOc13V9BErgCRADzWVikRyF3+X7iCC+J/ydCQC52B0FCh/BVmBitBssfDCcJ3DcJi79iADBhwFgpj2M29vH4m1iGw6B4+d9J4Q4tKEE3p+iHP5B5P+hHMphBMqiEvrmiR1lvCWkt9P7pSgFSvpSBfLFsXkC4XUi549oEZrdUf90D+lZJRZpAg40ctMTHsLyY9xHwg3oXNdnfRKwniZIXt4FxAsm4SnCG+Unf/KVQQJg6x+CflFKGUqmguAJX6RfggiYgvRlgujzvQBkwIU2vSgBAACu3ZiePiccPkBGIhbKIfLB/h+WgfJhouv/IctR/lxyveu7fhk+vhqm4EG4oMcDBPTVIubPhZObovrLSEOP/VH6tZhdqulT36A54+wXRQG+HNiYG0rQBxpWYRZiYfl9H/hrPd73Our+4SeOwfhlQv8B4p/Af8smDfxXjaDBSQm9CJzkUOCxhwnL/Zs0xQ+bf5wOevz4r8HBWixAmjw50ALKlQdFimQJ8+TLmAf/v/wDQjNavYNraPoE2e6fqJ8DTfnESTQA0YHSlrKM5BGO039u7kz1qOCqwAJEmZgKpS0RkAcgEy5DOUkAoGICABybxHBgwoNzB569OHCSxYtzJ90l+M/iX4EJAdxhwKnj1TJaaXYR+Niky8YfJRzcedIDSgACvbxg2ZPySRcgfYheucyRQABKT7sGOVMqSG9LYbhxjepfbo9KpnI9aO0klzvK/kU8OGliQeUmAQBguLBvXYnQBZ6dKNCixePHz57tHvigAAu8Nv5bxHLmwCX/GP9j8hpkApSTXcP/F5wmK5NFaIbGrF58Bx3wEyek/eTIMkAIIKBrv32Uxj+ANDhQ/4BIUdhYLJWMsMxxNHlxVjkgQocJRXFNB9JgHloH0orGgQTAIQNpphV7/whwSTEYVshjgI0xoQJl/X2EwI4CQiVacSbVk8pADBqJkgx1eBTNP41Y6SRlUtUHkhY3hmRSKB8J4ZGPJ8l40hT/lDTWQOCxiNcye4V3F0STANBWW87deRJZH9U5UTXJtfjPAy7OBcAbH2xzGgg0MfAal1rdB+RH01xlGZQNKtUaUap9dOVHZmpqkioeATLha1PKxhIeoXm020BZwWZSIh+haZIaJfChZqGGCmaXh9WUU4IMF90FIkJ3Osegc87OSehAhv41mLTheRTXQJwBkEuRjZUkEP8e/7Bq0gSuSUrZEzseSCupNCE5ELs/PeAIg3EINKq7HnnrLgxnsOQlSlmZo1Ul/3RgqUcAjMDHhdIO5l1EKlDCx0delOMXQiAmi5edgnphEEgigvzPtnh9ZLLCAgkgQAAt75LLQB809sWTJ5lLGWZginbBfQI5OlVTAl04gWIrqTeAvivh8A80AsnLksNx9ISu0vTtPFCoA72a70G2EmH1QBH+k6nBKKUqkAoyBAltYA5dTBZZDs1gyQgVwQlStsj11SFLeH55EFSRRNJI4YRnA0g2cSweRxqM0yJHYlO5FzaP+pYimUDXVP6RUa5B/Q/oJn3aEtbpuUvDTGND6BT/2DsybZLQmfq0Qyy9KvmwtWuOYEguI4R8kJ8mQeTaMZhMZHxczq5ss0CRpIqCHI2p9IZPPVylM+eZN9CkR2jSmHn2r23wj2lLoSCQmI2x2nWZ2p/OEq64UjbrQLC79kYPgZSDu3YfPVCOQBjCEJaYgXFElB2WcCdaL2IJADuTnbPELYIvulOeBNADLjSmRDRJ2hfEtZT2ce5SAonCSsi3PQE5jSjNE43W3ncQ0bFkdT9xXXzm85ppXAkAxhjBDjxSHNwp4zuBiAUBg1EOEU3wQ8EjipyEt5K2nSVkDMLEIShwinZ9pAT/KBYMY0IERIgQhmM0CbgEAgOOmOcqLhNN/wtPgzaBkHAqSTOJUuC1FDTZUFMvuddBEIaSRuwiEMZIokdwIjzhGcMQwDCEQAz1gGpV6yAL9AIUaUKWtsUEYwrrASFowkUuwkR6A8GZ1WbxD0h8EX7/0AEBfDMQoxEFfW08zQudgkcJveZ+JhEcDYmyx1V+BA6NAEEPVFAONc2pbRZ5gBp6Z4lATMGSgbkLAt2WomyiZJKBQeb/QII7QyUEeBbwRASEuRTxccAjBDAVOjN3Gg4cyAUohCG5pmKzOJ7mngPJpeXQyTWB0MInughAD3t1SSAOhAoxg5Z2LobNR1oLALsAQDnIMpi9rMghDxQIw4zxwyYu8VqXrEs1Av/xCyNBKiZDeadLYSJPmtxmlSywyvsC1Bp/itBWLwWJHca1C9v9Q0k4URPuDjKFGTgyEAPx30E0GR6LFCMA1ZDgnIpjkf41VSBKNcQIHnDUwEwhFiMQSBC3Oqdt7SKlPXXfR8TXVn2hciUEItA/giTMz4QNCygJgE7j2r46UikQLLgQUi50VIvwwZEJ9B9Un/pUZTxgCpNVg5rIgpSEToF3waACr/4XiBlQYSCSNSuMSiaAgf7EZz/xwyr3E1cM2dWuVmtfGjlXpZiU0aUxM6X0SPmPX3hCBWFNKFbv2ooEQjYmhlJGEif7j0Tg1VoG/Eev1HCQXCjTutmZQjDQQAX/r16LuxdVUkSc4wt+7pYmppyKmeAKE1ag7x+xEAgTLnDG2g7kBMaKT2RuGtsATyVTvPgH2Fw3s4EsIAq3M4nDLNKKsh4krFn11WZHYMgHAPABI6BbLrC7l73w6qLJTC4a/kGFIEh4CnwoK4f/YYgqDIEKweAuSJbonF34EV8msVEXhfkqn7CCBiUUiI8rt14Bg4rHpJqpaAgnzFf8478wsUwJKJGLXBgDBdkAxz82d6kFWNcihkWJAXslMmkBcAoRLhSJd8AwAhayUB7laiCqMQXvwlggjpzBDw0YjDwb0BBUAIYk/hFoNEtU0f8wHgh2/M+D9Je1MIHUXGvhXsqI/4QVZ1DXPzwNYIGc4CfX+8ceVjKOgWhAyV+85SojY4KltMKya8oyL4gQBV88YwSK9pLwzjqQGZQ1mUMlb0fJktRgGEKak/VuZ/8BjP0JBM58DoYvirGLGgukCgLJgCGSCuMT884Q4JXELZogiSowWmQM2UEgIJ1klHAAUho0pU3QaTaQOIBUPnoQq0/yRpfWL5UDuTdrOlU1UnUh1lOpmECwi9R/qAEnAbvJjQeS36cCocVJ7DAahA3nEbSis4a+RSx2kEyG8VnYgQjEMwYSDGAYwADAQPSJbf4PNJwYGLf4RxMaCZJYtIKpWAXZG+YblTV8QyBr8IWS0eOTU9Okpf8/IRhM4v0PlaySn8MEE9ZXNhB9NmYOvPz3UngBLoh7BLtq0EKvEFtsiUqYzmPuQS6qEAiGcVsgaPiujIdw6H8YQ5rGCEYn9sz3f3Bb5zU3d7r3fhA0ACMLVxhIIYZQhbLirsbfhmI51HC9XQjAFwEgPQp88dPXqILIHpFyPH9ygVV2Ld8gKbVH1qipe0hluqAKskASbPbgO/0gLZhAgSUuEDTnebNqcpjFRzoDyoZnssb4xzMWP5AqKHu0TRAIGMAwhLwv9iQ6H8Ll/6AIMhy6CozNec3/8I8+DMQW6V7xDHIRBER/tU2ByUEgGMIsu/APSuBHX6dBJgECWmckBxj/fCYBfAJxCei0Y7OTdQJhDVwHJVxRAE7WgPExAQMwCzGDfAOBXQyjBtg1BRSXZh8xBYRwC+cmCe2HBoH3B2RgeZhHfuD1D4AnEE3Qc4E3EGhgAP9QeQchf+hGBS0XC7nQCSmQAvrXTIWiBjOgBnIyCSGFAuTSdETBBSsFEhaggDRhJl/3E6vGOWjygBEoLmH4UpzRCL7XgXF4ZP9gLi3ABXwAcWimBi2mJm3HEicnhcZQBe7QBOIADFRgAJKQbj1nhE0wBIqHBlUQiZFYBTUHeN0nEH3QB7fwB0NwYpEIDJf4Ed3wD2PQcyc2WjVXc4hGd4UyArx2YcHwDKMWIAFX/2kgkYD/RltfBIfxwYH/MAcwAWkewSDW0ItEwRmiwmRx+BFsSCG8wAszoAInmHxpMxAjgF0VZ1rbFgxMxW3nhm4+eBIhgG6KKAnqp36S0ASY6BEhIH+SQAWIqIiMKBD0GAJjEAO6QA41B15OeBC8dhBqEAyUIBA1Rg66wGOh0QCY9kUzQYYfIYIsYYYNMhmj5hO8pxUtQCF4QBulsxTJqDS3ZSXHSCEkKRoT4Fq84DvTqHb11StkdRBe4jAvGBM2eBDsaITyp5Px9w/u4HPpiIn0KBAh8A/3uAAxEANjIBCjJQ/594/cpVQOVwXigAHosCWRNoI/sU40kWq08pArIf912jMTFlk5AwBqruENWrgUwMMZJikgEgACkeCWp2EZriYgOEMJLCkQDod8M9AJgTYQjpBn/zACLzcQ8PcTyXAQpLiY3TAK/7AAYvYR8SAQdHASjPAPyTAEQ0AGTTCEA9F+AtEJuVBgGcB0XgcmCsmQROE5PmE+ooBDpsOMV8M5wDUV6HAQNhIkthgfIuR8PvGLPjEkPTULzHAILVZnHvEMQaJs+pdQwfUPm9CTY2CTPzEG0ukR4KALUmEHPLAA3eAO3aCUAqGYJiGZ/6AIvTAQKTBao5V8I8B5BlBgx4cCYyAEu7AAPFAfDdApRLGVWmGAp2E+s0mgbgISc/mbBSr/GtsAjZbwDxE5EMbgXaNFCa2gJtr4D0ADEvRIAithB6nnEbggot3JAzxgB7rwoWMwDl35D3TQoZfxEWMAjygGY8EwA/lXaAbwimUVDNr3DxQQAqn3El+paZwzkf9wpKdBpO5CZR4JEiH1DzT0CE5hKG/xE2dpJJHQGgLAQVeBdbt1gHJADjqAAbzABcDgoP/wSeQWM4fXfjhRHCbkEQgJEjjpFLjwD3jqE2AwEOAgo5EXj/EIDE5IkHxXcxhAp0tqNQwooOOwiyV5EMEZYO70D3P4DyDkEQ94NGp2Mj8xnAPxGPtGE6pEEyAZHwwXH6FRXx5xC0NwiO5Ze+N5EHQ6/y5LoQt6qqd56hEgGhO6wANYkG4LNRBBkAEp4JQF1gQLAAf5gmmkIxA5IDaj+m/tkKRfhIEwERSNgaofkXEq4CgceRVrMCFI0aU00V8H4XoDAQ8wYVOyeRABcEc7sq0/oZEH0V60YEJqFwiMsoND6J5/qYcwcaIoAaIFOxC8ehB6eq0DwQNpMGqHiKMDMYTykAHywAtokALbwFZj5AjOiqkwITQWkKCnwQBeGHzntBILi60YIkoCQYEeQaoggQWwdRLKADz/0BP1oLJa4Vr/QKkwYZdfNFcH4Qc6UEKxoHaiNQQQIBCBN1oZUGA7YFmr2hgFq6d2cLUHi5C5uhKRCf8OQnCICxWPBpAFrxoEwTAClLANSEAUKPgTn9Q9O/KfL8Vw77CMNAEH/hQT2boSmnoQjzGvINGyymgPmvMTXuIIyoAdrtGkH9Gzm+OuSzYQizMQ+bEUsfkPgQsT+WayA5ENUYC0HsUHlhAEBoAMpLCDwFBzTviIPrRuV2GwAoGwunoQNGsSY/ALPycQOFpzBhAEKVZoLZYLawsTylBxavcPkbCz/8BXmrJODNBewtQFIuAKV7G8U+EHfisQpdAFotoYZBkTqiUQWsBNJzFTGmok/Wl2vxAFeFhWIyCEwPsPKQABEFAIVPCETXB5u/a6H3GrWHsQAPwPAizAovELMeD/DjbolL0Lj0HgwIWGtp2wDWSyFL2it1/kWnPZkMIkqY0bfAnqvfrSFIraGBMwtMXQvhDHO6RrAIV2EBmQAVkgEFeAu4FwC8+wAN35U7OLCwWsKeAADkpgiFVgAI8Ytr+LxBA8Ap0gS1tDE0qhwTAxkcPgLlKXcTIhICQMJR6MdDFhtEsBrVNxb8GkoKLRAChsCGpgBf/gly0MDKUrsYgIw9xGBgsAxOAQA3iqx3PKClirC32MC3/sx4AsyCYxux+Ren1sB78gDuIwBGKAYjWXfw6cxJaAtnywDT65So+KIRA6EHqlX3EVGZhjEiLZViAZm6WwrprrGmFVOVxRsv+w/1IrtQa/EAh8YAVr7JeWgIhLSaO8O1qbKRC6QKcFTLM9rMexO8DJzLWILBDInKcGCwc84JM2fBCTTMmUXEAixwma3FbwdRqnFpZxaAWWShnpQBP1xRjn+k4l4smkUr5hM8v/4C2CIBCBkAtWUFYzQAm+K6y7+w8RexK2G8AHa9CyG8h9fNDP/A+sQKupxwPDjA1YS7NI4AQ0GtABnc0P/Ip8wAlb4KSVUcZXkUWRO9IggTmi4MGrpCMncQmKNh/7Bg8h3CCurCk0cMUHwQD8cs+5sAS63An+7J7+HASraBK0WtDOHM0Hm8xRMbBLLbsf0cMH8ZgC8ZkPvNG/i418oP8NWJNwAmEFWoC8/IYhp5bTH0HQMTGgDcjKH4GlJ+0TLaO+r9G9PtGuMHEJFvAEr8jG/TwQb3wQq+iUGT0Q2ODMgpzQg6zYid3MIcrYf8ywKzGEWe3AvsMwq4CzqEkqA/cPfKtFovEbYdmyVOwa2Uqt8NRWXUDKILEflAbXgoUSzTPXjBsTKGAV7MwSKzmFncALaZqmaBAEaUrYPhHIzIy1x13c0dzYINHDgJzUgQ3Hk53NKRYEy7aHmM1jX00ZaX0Q1YraJwF1NDHOAkIgGnAA3m3SPUV1zDiv6doYT8KbqzS3A/EGboCc/NzCzfmXZSXQGI3RNXfRDf0PCFnI/7v/x1eb2At9EtDMEm/suw9eupTcjSK3CuEQUA1CwSGU3iYR3mDpE0TJZG651kgK11YzuPFR0k5xXgKhFEgRz+4Sezp9EFjgR8bQZga0zX/dCbDqEb0sEEbNEoE84AptB0Su0IiN2Frh4EVdusAbDGogcnMQDuDcIKw3ECyK3vHxCEwlELdxAe+8ElHsEZ5d4pRjJFz0S0ux0gLBqCxxWVlyEJ8qGusdHz3ABwa0xFRQVofHEkUNbX4OE7m6w0Z+osc9wEfO3QLBtB/xmRIb4RBuAF4F5RcQjFZzb0earVl+GugTJNfjRfExW/9AICwK1+fq2o2hSqLEBCcOQ3jlIgJC/+dr/rYDwVR4aEC2nooescB/DW0e0ejMTdAoOsypJ+wDjpA7jBL+/A+N/uDL/ugRbglowGtpmw43QCFb2Zq6YOVIiuUCQebMiA+iLhDnXeIHsQsfOxCXQEMPON8xAcoiITQ/4QBr3rnopAF0vhKnfhBQhwg0AAIqEAt8AK0QFwyTvOwDEQ4/qvAU8KOSQAGNLA5TqbrAcAQCwpgmweMHAenPvs1TaAnpgAP+sBJxOxW2KUxgXu5Kg9vqvuGZluYwwXCyrhVAILKvoQEaMA4aUArc659sPhAHeAkJaHdlVYKtMNjLXgWj8AhL/wjT8Aj2sPTvcApSIAwrgAGu4ApmQP8GF02UtuAuGe/sG++7eo6NI8ALIB/RFDIL7Q6gwpTiKPHtcH3XAoHbSD0VVPsPwxi0NEHT+jEQAuhgI7sUN3/zVJfhMNHFArE4teDvL2AMuRDGr8hIM5d9m4Cnj6Cnl+IP53AOeuD5/+D5eiAMNvAPXt+DU7EN4nAQTmvVR8/oz/7gvPyKUzgLskANDRK9cRXjKd8YONT3HnHq6JvZAxHLba8VMu9EKIGRM2ENNsMCxmK7mKMBPpDzVPfFMdHmAiEHKFALePAGd+A7EveKLty0NLcFUyoQ6P/5JkEPMUGUOFmd/xAOmbACmVADWwALGLACK6D1ADEE2D+CQQge/Gf/wNK/IAaAGWgYEc2IEWpmbJv3LwJCjh09fgQZ8t84kSVNftxzUiXHdv9aklwZU+ZMmgTfdBxT82ODBqp0/vQIpKMEkA3+1eP45QtBVgSb/BOlQapUUaJK/dNB0KjHEkwudOTwjwMDOSho4HkRy9CSfxRnGOgITJyUb/8e+UOo5yA9j01uAQUJC8fDghwNJnxoycDiiMHUWFETbJssD4A7duBIwPJmziCHdQYZALRJBx6Z/JMR8ibCsGJjpiZozahRn6N/LmX7j6jHrQQFdEz1b2vUqOOmllIgaE1IGacJtv7H5t8iDgNQ4HkTK9cIKxVHdEpI0CFBcRXs/jAvkt4p/00r/8akN4jMwIEdDT5siB+igU4zplTMBZphKqPJApEG+AdB2xYEqT2VQkGAwZnmYLCHVkra4SAWDqKOJhYuieMgX2yDbrTlSgrunxWqmooqUWRJQJysSvqKIFNsNKW6M0BQIZcLl3BrIY/megcvk075B4mDQngqpPdWqsEVMqg4aCC4DIJrMS21VGwiNSriZY5hFEDRNAnPRCilGmPqzSMf0EQoBzj/6eIkGFQAqYXnapJBqH/QkXCRORHSAgg5U9TkBg+6SIDRBB6FUBxyTuSqI1Nu5ODSAaIAIZZENhxhhu94+YdUjij4oZmD9NKLHr4wEOYjcDrT659BxKlPyP+Drkxov8UUe0jUL5fIoAsNyFTpAmWZOA2PQUFLzblKZmpTuo9aEqnNmSyQEzAANoNtQT4ICmAXTP4591kGHyBoKeGgimqqdjQQRRtechHnF5FK4MgUNi5dZIAzojikFRZmWGKGt1LgSByCMHCmVpEesesgSFLszBUzEMqSoyy31BKYICj6cgZtojrJkwL+qeSCPZT9iAh1+eQIhn9KU0lbjt5ESIOSdFZpim47w8KjBACbBTBl0KWJwpM4kRBogrQ4qIFwrJpqHg2GeYVUPsSpYtaD7CCI33/K+Aezfy5lgwNOOOCih0Ny+UfhUMGDqz4DGL6CHYJs6IgHgtLzSPD/n+pKkiN3OKovPIIeemhLcSwheYRWVvkMJEoJKkBZl5UlChCtCOrAD4JM9wiEf3Bg80yzfwbtXG+W+2FmkAhB0xRB/9FzpqUM1KlOk9IATWqOjGJRgwOoWoWSf1rJJREs1jCeIAYY4ICDtt/mghdSFRa1FV5SWIxhRlQyHCQkgaK09vT/ef+f8/8ZqCGQHRrZO0vSKYVnj5AiCC7O0LmWvWwPEviC6Oxgh1nJAUETQAghMHYQN9iuI1+5QLg4c4B/cFA1tilH2mqCC4Sg4CRretqeZlIEdwHFAcJTV/X+IQ3hUABrGvBBVBzACecRhA+8cAccOpIb62FPe0e0V91K/6AwPhjAVBKK32iiKAmHhMyJwKCIFWZACYdRQHNascMZcnGBlrXsAiww4RiM8YxAEGAAClIbQrYCPAseBIX/0IZtOOizknzrJKIRzYI24hEXiOQJJTkEQhZxo5qcq4UrOdo/XiGTBkTjH4jryCFzZhKkOCBePpBKF7ZBkE74yBC8wIIQ/9EDfhHxH7MwYtvYwAku8IEPM1hiKyyRgiNwZJAI+eVMdAGSKB6kCTbYwj828Y/lUCxW8PsIxsBQiIdQcTHAAIawZrCPjPivI/XgSQPs8AICXiAXe6iEDLQTix30wA0O+wfqDnIHrQCKjnW0I+dOQkOPbAAaIeHjZgKJT/+EyACFT9jQQVQ3kzcUASRCSRdB7kk6zrjhW8XYhQCykQYlaPIfh3yCzX4yCYQ8whVYK44GXrEPgjivFeD5RxX+dJAloK0MF+ACF4zIAG0kbQa3VJiQANcRfWmEIO+LATQPYsmZFPOoBFkfQSj2D2cUTnBXxcZThiAJ8mnJS3yYRTpEIcmOUI96PPmGDghYiUo8gRKW4MMUVPCfD6BOnryjJ0FSsVCQePB4aJrkQbz5kYRugKAgAYBHz/SVlIAmQx1xDppKdC5MvOENIBBAIJ6QErrpJER+PIjo/uEKB5SCXlI5wCu48I8ewjQXzgtEFP5hszLU9gITuN4stLePC9z/8pa6zABBkppUXwZOJPag2FRr4tRp/IOpSYgqR/zRFDsYbgjl21t/LMKLV6DseDwBJ08egYICoPMClGgBLygCJIskggu9i6fpIAgUGVomsINFCBAeq667qsSP/zxsgC2DiR1UdgcseALMWEaQpfVXtiEJAEk7YskueHIcoNTAPObAC10h5AK82EcsSlCCMpBYBhMYABdmwQYu5OKnPxUfw0ASTIRc9SPvkKozjUsTHiTBLsr18QQDZ929GUAghqBILFZRlVd48azhhPI0yEvGFrTgYKHqjhYpMYsWrLYmxuHNSrRXE2xhS8D9NckOQCvgzhhoNSBBs05iQVnL7uDA/2Qk4x7GmBo8nWQNJ5LwQUJEwgrHSyrziAc/DEA3mBKks14bcYlbMAEucGAWT/jtDNDwRITE4JdOfSpC+HIQ5RLESNB8n+F44NSrpiKpz5wJMv5BvhSQT1Qj4EUCNOAAV0DZ1+GkQQG8ZzfucGcGFtnyP7ysoDh7hIMw+cfKZuICRs4Eh2z2yG+wLZMd9Pkf3p7JFP6xlDdLaM5vIPAb7MwCPCdiFrx4QizATZBEcgQOcDiRaP8RaKhK0gQ3PPQqkDEEKv0DpuC5UCsowYtK8KEEfmgBB3jh2xdz+iPE7QjGEUI4qXZkfenjwayQZOODgDqATCUIrEtC671RYgZaHP9COuJxgyc34B5QXsMYCHCI9b4cYS93Cy9WywCdjCO1/+isuvy6bd/YZhn/ePrMrCUTcUe0JjA0ybksq+47twzE2tAGF+4QCy5YC74cIV6IGnEQfiOku6adyjBAsYp/8IPDCGlF3ltxS9aidxazmEEsXiw+lhIkD532iMaL2xHl2qMjpxacP1JxVVWjWiQkrNhJZF1k8lFhBizgAz9ecQM48IR6N2+ALshRBWOMgAVY/nnCQoXrnBLdy/E9w0f4KIoD9N7opWksQTZ3FDThl+nq2t1PeheWSyXrIEwQt01KcvaPmMAk1fiHMgps5xJ8rhKzYIayZ7EKbUCNCxOYABH/1BYJ0cUhDXGIw9r/4YWDrPkfcyj0J+MxP37YnQoI95FWmIHTKAMmaAGXG4ElmoFWYJgMCC7Eq6qiIohgUrxR2DhSyzyO4IHJ48CSgx/FOwkSwrGTMALxqLUUQIMZ+AdD0AYciAbTW4NfaKNYeD1R+TmFkb1QOaVtIADWUTaOUAKQIIl2OAAfWJ6ju6OqGR2PGKaDGD7bKKRn+Y0pBIwicCiRiJCDUJCfMAXDWolpOQhv24GJKglUSADrI4guQEOVKAIL2IESMK9KaIE8Krx/YAZoWAUW8wM/6AA3EIBIaAT3gz/5oz+ECBE5IIhXKC2425p4uIKD4Icj4LBS6gSY/9oiXnA58JmBU3rAgygEgliAf5CCj6iqqjIJzHuER8A8y/uHyQscvMCLpCK5kFgDbFjFkpAEgjjBFKCCuyEAcNAFHQgDY9gOG5w98EkYu+kEEMuAIcCCoTMJBJAF1FIeI1Qe1ZI2y3jCzYhCOFkabaNCzhAKZzk+gvgKJlCDgyg3j8CMCgoJE8C6j6gGy0IXN+y+SkAnStAGZsgAEOMF+NqHv7sXAQiARgAE+AOERhAAL2DISXBIgvAFOUiAOTCBVygFRqwKUPgHWYMACNjIfnQeW1oIPhA8G2TAIejEfxiCjQwJU9Q4EFQJSBCbViSI2oGfCEgfcFi1nVw1hMCGdf9IghhAnPT5g1+ASY6otb2xhGBAOl5AMreQvRsEn9lbuAxIgQzgh3BQgkr7B6KbhdvjCGeRheQ5QuUxAQShBE+4xXcRsKn7By9kEKEAx4O4wnIEiWqzQ0P6B85SCQNZmrbjiDU8icq6iTeMw1yYBW3YB6H7x8YkCEvIBe/Zjl2IhIJshAAAgEnwAs2chIKkATlQAAXIAxO4SA0wLVEQAbpDho6EgNVEBmTYhm0AMbh6MVE5JZ0wxVP0CCWpnaP8hwVYgD7ogxCwhZkwAjBQhIM4SlLoiKRMAUP4qX8AKk2kzhFQi1qzymbMAjIIRQSAJY4wndn4hwDAAwSwyP7BIeX/MUs/sIR9MAaCAKCZIB67pM9nIbqTSLqS+EqCmC/OOJc3xLNKKIBEYIaw44d9GILx8R5KSIRc6A+CiAXtaL0dqIZJyMzNLMhdAE0FeBQH8KRSeBEuIIRVWIUrWM02aE1k4AcI2AdLiAVbEsAZAA8ZS0mOKM6DOIF/iAFn2FHA+AOR+IQr+IQfRYhPMILk9IhPmImhOoghuMontYQFvJdQAZ8SoFJD2CUHvEotPQIs+AZNQIASOQgUMD04IE8ueDtQAqXlUSlmUDhCIB7xZMvDcsszaQEyFEeRuE/AqLR/WRtrcUeOsLrgI6jVMMwyYitKID8S/QcIOIIhmBxMpASS/wwVNVCDKbBUXMo7PhiBHQgAEBAHBViFRzEBE/DQF9oGFTCGKwCFK+jIVYAAurMEQ+iETc27WhuClWSYlVzJkiCu3KQxzjACI1DSjlDSTyCFYiUIZZUJMPgIJ82AWZ0B7wEqPuiEXeKFZtTWDMgCBywESWhCsRgLhLCOMiVP88Sa03yTDbulRHgGVfqH2iiGk6iNa/CFdTyJsRKJKITLmNgv//qHcIQTBCDY0ahT2xFMkJCtdPlPPvCcMvowbWBUglgFEuAHeeCwvFOYx7BUTPXY6BsBkczWApXYVQAFaNiGIcip/uPHFLAEyKSETqCEl+IDKshWXm1SjsgChMgJC/9C1k9QVqD9BDAAA6AlVqAlUst4wCeN1hddzFnbVgd0wCxAyQw4AjLQl61wm+y5HhQjU54w0/JUxC6oimFIh1CY2Z/6ofcc03Yhx5KQP45IqI/YI9uxupJ4JAmJkPvcwp+YOrx8ljqxvoQFCez7B3QjCINqmXNqKxbIBTqgA4IABY0kiFjlB2bghV4cgf/oWEtVA0e41ND9ki+xTj6gVUpYuNTFxNVFXZntBAPIAHkgCJRUCTIoiWDlDDuIgW5AUuUstRIMAR5Yy5nIVZX8h+Da0n3ohGCwBHmQ2m6dWm6d2iEoqjUQBOzJETa4Hi4oV7ANgC/Yhld4hXjQsFp6Ud//6oQWiIVdmM9/sLN2kQm+EsKAGo14dN+Z2IG3rc+PyJQbSb6ZKVV4WIlvMdw3mAKHVRYzugAYsIBcmAM6cJp/oDuCuII2+IdREoggCIZbmwJM/dwO9tzRVZi8Q11LUN23eqtcsAQQkwd+GCXZ3dmPeMAY9tUJrAls8AgRfIR3wIahutFuED5nsAFnVc5/wLwRLIkc7YiVRF6ptUpDOCXn7dYpzgKqzYJtIIdwst4wzZFF6FrriL9IiAQ8KE8InoVDgAGF6Q8BVDheSI1dQAg3JIjo64wDgDbbgSeQSBc4tgw8mTeQ6E+8NYn/7YgdqMsLWJkkDIlFgBqQSNhGRqy7/3U0lnEZhJKAHhCHeTi8g9jkRt1I2Z01hAgCKuCDYKCIKQgEznWLBXypa0Xhl3WifeglfmgDfvgHMaCJTg5FoxIuYKIqHeVlxsNhjkjFDCSIbwiBf+jdZP6HEYyBoVIEMLjRmFicnEUIGp5iq8wFKsBKeajibciAbeCHVcgFEIgDs6qDt1kERr4eBhgAFQAAAYjnQIjMVqgIKY3WBVzAheMDFZDkf9WJbCQI+q0Jff0IcXisDAFoCwKCP+aIPQUKiG6+g1gaGjkJ6YDkdzwIzQCJY1BHD0M6REYoFSCYUIDcf+hkyt3IQqDaf8jFXCSIXKSPf6ACKkADQ7jpTggCxf/I1tjdBo5ECFk7CAsWiV7liMiNCdzFCyTGYRwjIeVCRd7lCGegGBLCBnvAhuJUBEVgZpXIzZJ43iGA3iCITGaQhyMQZ14wBmOIggBIgzXggWfYKU5gAGaYhQGI0Oi5pf/YxF2qtVmVWT6ITF6QNyCwgDdbDTpGCC+sN5kwvs7QPvdd6ChotoNYaMDoMxXwE4/ozxs4ibxFCN2xkY54syuMhXB5nZIQU4TAmX+AR8CY2x4g6UPgBE6QuU1W6YPopQeEafJxnF6JnAYkCDF4TYTwyMq1YKFuA+LuJaAYRcSDSQz4TY8o5qc+iBHEhnBQ5n8Y2j4wYoTABVvkUVv8bpr/8BuPAGWCkN4skAfZDQJDUGFxIBVeSIQ1QoFAqILYjE1t2AbMvRfBCwZdytZZSwEnXQwHNIBgoO8L+YcrVB2FBmhBIWSZIGiZKCTv8ojGVmjLXokMAe2fqMuH1gn7O4gbYSSI5nDAoGsUJ4jWljOCOKQa2RCCyR42mIOM6AgSAAm48JiO6EShPojjBgkg9wij7oj5SbyO+GqPGOZiTq6KSUWK+YZ7IGYcK2apwrFhbuaSsN1OSyakLAnZ3e2/pgL4NoQSVuE0zwX4vtYBR8pdxM7MTd8C4IPIMlR1K4n8VInMWQk2WIQo7EaRELfLNonSPr5CtA1FromrAA1pM5AP/2AAf+EEBZCFeOgIIt9xmtBxjpA1Cz6CXkrvj+hWkaCxo9zlACK1qjZmjrByqbLqf9DydwjvUoP1kNiEaiYIMEjamDiCUP+H9tbSqG1h2ZUHcD5elVza7GRaYDilRNAQjsgQ+QWLf/gAPAUN6ZCOQA+Jzf4HOlLszhDo/f0IxdqMUz0JZ9c2kBDpHjiI62GbbUiAeUBqjiDqkNibmmhNlaBd4z2IUfKIYAVWJmf178bhJ3/ytXRqKE8uIyGh4UWIBciEkqhik+glUP8HGtbtW9b4XhKDnWVv9Ub2YL/KXD2leylkhLjsG2nkD1CXjF4JfGUQF5cJ3OIMFu+MdRYJnP+x3/ojCBAAANCSZITwKHd8mxypbTrQ5H/YdEznCCOH6d8GCSGvXI8UaqGeeH4X9Z0FhV3fiIDv0SXv5YPABVlv6vDechFs5igXwYZ/h+TK8lV0+AbB9X/ocp1VCVwWgyOQNaEm7oPAe52tYulVdshchaSJlgbv+ZOo60CVvpK4Y5Ow+Y6ocJnghKSxjJ2fGeZbCXI/CQ7YnXBPQzrRS48I+o5AgNUKC+xhAC74AE6I3An+h+ZGCN/+CB5XyavvCKknCKbniODqxBrtiFHE3YMIxQggrmRe6o64RYOH8sxTrqrGBopBYo449UERatnH5aEmiOY+gioOfOjFpit4BQb/cMcSyIEQFzBEDFPPP4lQCAlCD7BA7gwE2FOA3gF3iQWvmInVPgiAKPVvIMGCBv+5AVFQQLWDDrn848BAIgMEXO68CbSKDomByJD9yzLECMEhBQ0UTGGwjUEIDg2CJFiooEmD8kK+HBjhpbMY/3zmxIbr3aN/uPwZ/fcuaVFc/4oShEpw6TukSHMCzfkyi1aCR1iyJMgS5NiBbcSwFHNk7ZEsWTK8TQFs1RwTCAcyGVEQU1eDO/rmHAf4H4NFAzk41NB3B99/fw8aHizZYYHJOQFYJkzxXy6HbwjGMhj63xeFDhkQrPiyi6hX/+y+LNDhyUHMkxEzgBjrDe83CED9/+OH7AjNkn0z9HX5L6Zl5P9uOpTSNUbPnE6x6eRRcKnTpUWLLsWOPSl2p5lzctVK3KAYg/wIgiQLAVmbNsjEDGe7Nos8cVxWuWbCADIMVIIE5xX02WMIMliQYv948NKCKrwEUYMX/jNAX7YNZqFltA3EB4avDeTAQAmMOFksO1TT2xvizNERSIUgl0JNg2XBnHL/dATTcv+oJRl0L0nn0AJ9rdPXVf+IlyJBRwr50nDMwRecQ2DNN599bRzBzzZHZDDENgbhQOA/JfzDYWOAuXFhFwR98c+aBU1w2EQaCuSkZHrp2SdgdRr0maALgpaiiW/C5qdDda74xRsC/MPbDv+8cALKNmP+o5Jl7S1HSkEQdKTcjgWldx4NBp1AUFb/OKOVK+po9Z2TOxkkwj99/DOGQTMBtt6PDimH5T8QtKElffiJUcgQq+TxD4oEoQkDmphxONgdluX5jwMmdiXOP4ASBK6iXVGo5yX/3DBZted11hUfILYyGWrjMqhhm59R+4YKsYzAAi+reFmTSc4NRuVBJLgUlqK0/lRQqxgmQS+CBh806kHFQpAxscYiw08ezSZqEAss9LAmZrv801BBCPzjoTGEZvamZPNK3BefNWcIGKSZEQLzQL1d65lWNK+Gc4UGVYsmCyqoMII42/Bz4xAEW3aFoqUWJN1ODPu0ap//ZviJBIbMKcxSwhojozE/apNAhyyuvXQgQdXGqdUEGhqtJ8p5G71zZnP+s7djBoH4WU7iOjSHzHx3JfgSA+WgDAACEHIFwDOFyfhkYhvU6tZaUWCQrgV5rfnEv/6jsMars54xMm3H0+ziBckBWN2mM1j7IQ4JLjjuF0Lqd1cEYEjgX3h0BaiHF0bSJ/LI316QBbd7sE0oqyjw3u+TaU0Qw5aVjlWfQmRmMMVZtr7663PgUEUCcP8zO0FyLxT4S3Xijff2lqEMqe/noalBH9BTGgYCh3/EIQ4DIcQhdrc/BgWgeVohUA8GYwGD+G4EFVzgQDjxD8NwYhWrGIiyblQq/+1ZbCApXE5+/sErh2DNIJw7iHR88rCDyG8gN/xewwrCsAhQ5yXfq8A/oCTDIxnxIO1Bi8I8krphtQ5haEMbCVYhjr3Z6h/wGIhrXqEArQivKzd6YGbW1RcUEKRcAxkNggY4ogMesCBovBAM+pRDyUjQIAEETBH+gTyCfKaOBtLLZ6pQkEW4YCCGEcczCCEJMhTiUkPgjxhQaDXAnIVTLoRhV5BYJFb9g4cFgZX3QpmZrASxh6WUziefRJAxLGCG6SoIWNpTH4IQazlTdF3GpJixK4DiCsYQwC5sk0WCwC8nAeDbs8h4IRZkhggF+aNBpDmYNMAhmwRR4EDyOJD/Of9TK424ECH+UU7e/YONAymCAAjACQ+8EwEekCcCEECAXTQCEI0ohi+UQAgxrQJUq+gRsA7yka7E8CBiQ6LDJhOBCOywlEB0GFBu2LDPsXIgSSTIJo40w4GMcCVmyVKx0pa+XoIKVKCgwzYIgTJ8vcGBfaEfQZZZs2ZByDL608pO/aTOgVjAcNuLo0F6EAWDuHEwZnLIHL01kJ46yRs5WZpp/mHN2mXIqVqp4wbb+c54znMR9cwFPq0BCH1awxsCAMAOdhCIEeQiF7wQxxXokA864JUOoACFS1bYF664hSAfPYgoC5KMgYxOh977hWJ9qBWf7CRVGS0iZTm3gMTm6h//TiAIp+wDgbWlLbTom+LrVrqKKwxheV05p87spxWsflOoa5zM88IpMdhKpoC/g6ZBFIKCF9RsnOOkVx3T6Mcz/IMARLiBcpX7AQJ4whf5PGsjGhEJAQgAE24dQRWWtQq+5sSvLxnSc373sM8dBLKm7MsCOjqGwZqBEYWYEj/aUF/R4hd9VQTFKjjhrQHgoCDRy8kxDaLGzMwxjPwbCDUBs0XbSga3XZFwX4hKkKNaZoNdQWO79qdG4P7DDxb8B2//oWGChBUHCMBBKBBQhWeEwR1hIAQBcjEEeXgpY6vQxmlfgrBhiYViu5LMAib7j1YCJgT/sME/wsETykLJazth/6xBGGrZgZBvE0IYxUCO8JH7fPm+6OPvabeRiyigjHgi1upABnyQAjvENgrOyQvQ2GCCWKC4g5nzS1jWIDPyzZp+srBDCMHacw0kAOAkSNAeGAlvDqQHIK5ZgP+BAADjYBXIUNZMYtiemFwSlzmJj2RKRQJ2GISIehrsQCKGIcy+BAJ8DSjAjiDJIYhDHLkghDEibbij6g+qDHrBnf/BZzD+A9H/0DOEidmgoLFx0S8hgkxxBtxJu9am/9A2o+VYkFPhTKovOTDfcJAuLETCF1Ugg9UwNcZfzQfIUnoiftYiE4P4yjgQpmwpZSiZeFwhBYF4wy52QUxi4iEQPbgDw/81jDJAD4R4L1FAM/vC7W0f2yC+gFQANr6LQAzkEB5stqkIcuJ/XJBvkB7IGv5BaIdg2H+udVKvUwTpqmIQQ57oyw3SVYt/0OIfjUCBONjtwgwUgjhiEBVgMnYQe78QJzO5ib2LOFhVF2SjOKPGP7iu2SUfxB0DWUET0oVqkI6wCo8i+C5KE4U79CDuRvUj3SX+D6yymUEgP88ZNm5slBn8H3v3k91xN0cDj0jYBAFE84ZrGTRiuyC+cMjJJVNtgrBYMp74o3CFHimDRD4nWCCIACav07sXhJv/AMQ3q/A0EQZHtBbTmLyN9Q/iEMctuj+CPNpSiCz4HhnJcLLWcVf/g4HA4h+wWAHYXLiemXj5H1abvkfsG58rkGAbVfBF21/w9oXHPQpRwMMu8LDzrggvFJaxafNWXhA2K5tegq5ZzQki7d+533YDQe5LUDZ5DGdGUh0EhWnF6A1E57Hez/yDaeDBH4GbMpneP/jC4SnKGzwDAYgDP3zXHOhVRyAMCVwBaU2Jl32JPERSJDkBGeAAGZhBOITDCqzAKDgZBlwWhhxfXxzf8SWfQQyC8sHCIAxC9fxeW+iHWtwHl2wJfZTUfFxB2vAXIYifMfSAJ0xhFATC3kSBIXXF5D3gZETQP7SfZcSfxAhggxQbCJDfQJzLGOIONyjKxalhQZDbYHxA/+iEnuYpW3U53smcR+nZ30Ac1R1iCHYVRBXcwNNswxVcCg5cSiRdyhVA4hUwwip4wA2EwxZkAhJIgTOcQzM4gzNUQDOcQwVUgA04weiIDatNxg3mBCtqBSzAgiuIwKX0Xu8dgVqoBZcMRxKSVJaI1nehFq8p3D+MH/KcAWs5xORdQgB0oUMgQJsYBBwehAMRwO6gAPKwoaJIEzIyCLiFzr4dhDTAASvkRAMQhDk6xB+hwCU4Xl8AoLHlxAAJIM7lnUN8Yxx63urh40BQYLI9gz0aQz9eguDsHf/l1EuIW0EwXiRo25x9ADKewSX4wkR2nKIJwj+sQCZWgBScQ+f8w/8o0kMNrMDyZR1i/cMmNNlguKJD1EDy7WAOFsQO/sMg/KArhEMVbAMyAMwITgl9fJlnLaHsZYnlACMOEAI5EEQdFMQ9GkSDRchg4IE0akVSRaDRECDfGGTeiGNOrIE5emVXgFsCDkQxnNFAVCVSEcQA9WNBbJZWIKVl/NzPvcT51dS5ZOU/3KVBMKXqdRNBPJpWcOM/1IIvSGQAKAEFZMI/fJQnghIR1UAPDgRkgk0/EIQIOIEZuALyaQVM/kMOJkESCIMeSEbyQWYsuoIS7AL/iQMjipAIiBAyNGETelZ+0SYEhCBR6tUsigMWCGAdGkQ29sUd5l9TgmNxngcGAEb/A3ylVvzcJViDQeyTZARdMxIEISQVCszRO/5DpR2EAfbl4llDI3hDHgWAsgXdQGAAFiCnViAaCCgBzvWFNRSQ6vFlJFiX553nS5yLXPoCM2IBU3YkKHWkqq3AQbhCDw6C182kZhqETBJEDdQAPaxDMzTDDxREM7xESC4oLCrfTFLDaV4CclXBc52TE1hPKIiAAuRBAuTBHLQof+UBKOQBs6zUXsmoCG3DELzYLnwhQVCAGxlSP96fQwzYfRpnZgAngiSpn3inVijnORLENfxDQvYFWebE3lBZAeIlQQiikwSAlRYaQTzgWXYpQczSQEgpX3ZFNvyDEgyEUobBP+wc/yIMhFz+HApQAAakog515CjeYIESBBAmaD8AYUwexA4mXw0kgR6EYoU2FmBQqDC4WoECITVgAHXmhJ+RwfZNJAr4Ag1MIPd9nOCBwN6hQCBQ0z/+A3Kyqp+0o+mAqVZw50u46bjMEQicAXyazpOiY5Q6BJUeYF8ohFyK3kDEKUGcARo16WAM50uwaXf+w7IWBMgB1+A5RGYOhA4chOq5n5TWal4iQi3QaUEoQRi4QiYORDOEooYexCC4wrsmAaAC6kvAQhLQQwWcww9g6D9YqL6yCkRZKKv0K78SBIb+QCeSYkgm3w1cZHUORrr8EbE250GYhhIUW7QOhLSiJ4MM1/+r/sOxjstZNghyTV4tXJxUWkbFHqlYDgTrRYNDeOxkKKXExEHMoizh5YSavoQOrCX50GlcEoQSYCcGuIIw/IO60sO8YuRAUMMKTOjRfiS7Li0sRiiFiuIPtMrD7KtBBCzXEqzAskpHOoO6rgAGaGtBaOw/kAFgVCWmHkQYYAHI1qpBgGyf1O2RulbJ/uaFgJybuqnb8k2vFoSUAoY+aQVhDsZFnm221oyUuuHiEkTDEkQxxOUlLC7kWkYCdQWdui0tqEKdSuAu8KwOKEE4JME6VEASZMIKQGjSziSjYmif/oOqVUBISii+7qvYbu1HnofuNlYzJIErmK1JOoRWnan/t/ycNBbDA6LRWhqrouzCz3XeYOitQ6hqX/hCrGLI4oJpMZBlMSwpYAweGg1pzQguy/2DbqVvQbRc6unsPwAu0OWE5LqKZbBsPg7G3P5DrNKA856HAt0v6B6EJmgFdqKAEqwAPTAqo5IiRmYChm7t7hJEq0Sw2IJSn1DwOXRkOFCAEJxKF9IvQWCrZLjtz43OzBLEHMVqCANGHhLEc+JtZpClyF4IDTNOr65B+xqE+v6DDjPI5+JOANvW+8bBNXwuEGuFNYAbDeiADmRkaHbmP2SCqrVKRyJZX1jUS1jwo1axQwToKK4D61LAFtCA9nbFmR6EXJbnP+iA28KaQXhv/4PsQn7qI2DQ8ZHGqk295YWgkQ0PxhY0yFee78t1hVjGb59cMUFUl0Ow7PvmBAwXxAlQWapkBl/ysG6pHgyP60GA6afqQDhkQib04L0eBIYm8kAE6AU7RBZ/JCsXRCpPMO+C4urqQdnSALAeBFMiyCGn8EBkw7MCxilnBpuasTMRKy0QM7GOCLj5cV8k5kFsAQEbhIUJ7vk6ySYritIOhHQEXbNaBvf+AzocBA1gM4LoFg8PBhL/wy/4ghCYgRP0A9cZ7T8kiUGkctYOBNbZM0EQESxrhT9DbSpb8ewKA+ueQ2KSzz8kdC4XhDY7XjHk589JMoIUAzEPBiWDrjXcMf9g4DK9YHRmxGxXqHNO8LJlELAgaIImlLNDLOeIqMJGx7BkZMNwvTRB0Gn45gQ2FYRuWRg6XAMkOIQCpcI/qAIg/II4iADYOFlBVEA9dwURQfVLYF0/Q+1k4HOqVYBICsM51LNcCoEQ6C9zasVK58RCD4Tnsmk2PKdZDwZMWwYkK4oQfLTRpMJQSwbmIog0O0QOG0RL94U1OwRQy29Ma8Unsd44oYMqjLQyE8Qz94X68rRWCPZAKFAcjIITsMMfMJlBJEmS0G5XzNAM6bM+P/VkkOIgrEADAyqV4bVDAPI/qDXMBt0JMLZWaOvZ/vJMtylgfHCDwLVkaMJkGwQwOwT/WQ/Gb4t0Ao50lg5ESUsG+bA1QRCyIP8DYLOvVqRBKoglIjB3MEfASI9IAnITUVm3s6JDNqCD5w4EIqhCBACuXjsEHAHGNYgzJEQAN4hjN2jWH/zBP5hBCHRDxLjaZCSJaL6EU3uxR0Y1YKxDEgyCq61DJujyQKiiQSACOtwv6yXgAzIWlbn1kRj3WNs0cxcxZRO1mFJyqhDuZr72DSamXeeNOCuyZcD4S9R2g0Q3QaCzD0Npeb8EjxNETWfG5zL3Qs9zZsj4dQ/GitN3NtAxeBsESqZeQcg3IReEG/5DKvDAGoQAO5iBLQyEItiAGei3Vnw2aacagkvGVPMzg78u/0EkwVKfR5IPd0Fk6SbP9T/kuWW4tVhyg3D70Ion7j9oQpHUuGSwcCH/g6D/ryr89HpfyKEf2aQLs1YA+YUcMZSPtaYrJoPIODp/5cvmRCrEgU+Hs2CnAqAjiHwbRMvFUQHZARxsgRMoQkHw95gPRDdEKEEcOT1LBurWs6qJplM7tWgSkYEThJrnM1PHaw14dpK4whYgQmH1hTirnpQSd5CrwvvuOaYjEGULtUMwDDlqRaJDDHxXuxEL8WRIqVvriZH1dUFQt6Jwgy7EAS6kAbnnRLfnBHoZRFH/A5brODpL9z+wgpYXBFCLs13HwefWOLXnhJVTefrCgU6vQSbQev9BgLktaDbYmMEKDDhB0MM/HDmaP7UwKDuDkHaSaHOTrUCq8HtBGO0MSTpBCLddq0IqQPyiZ8ZkA/VQg8NLQMK4qrpW6LWUD4Qu1AyMM3pmSAPOPNTX7ny8+3WKKH2+SwM5skIa2IFW1HV217xiubKJE0TQr+/Zv8TTG4Rdsx43ODxBhD1gvOylD8TLxlEDLAAY1LpB9HfHU4OSlblDhLGS/UPIM7XMw/k6rIOxp1pp+/pA1LPiJ8nIQ/5A1IArEHClk3aNo0OpZ/nnx31BhP55TLbSK71BCPYpDAQPpALBg7bp0HlXfE8anL6fiDphDUTRoy+QVz2DtO8BmT4c2EH/NHQ9QWhHwkeAdgi8XWttVcO9YCs9N3Q+OKheGrj+NOsCOiu96rGe2Rs8K6i+ZKge3RNEDnP5ZhG+xjOZGWRC4B+EfneDEyQDKSSDInTDApyuVkD46QoDQFT490/Yv3UDESb8J3Agw4QFkxBcd1BhkhrUzETgweMfR4UfQX4E949VyAgDYyD0GJKlwlQIRw4cqetfHIWnBr5s2dLZTlU7FyaU8hFSqlRpWp5AeFKhtJIDcbGEBJRqQn8InypsoPXf1q1VQ35VGO2fNDhw/qH9hzQnzqkcWUlT+IPpj392Q9r8qLbl1jUD16RRK3dtzYG6dLEiG/VfhB/O6NqdmpNm/0LBQBvEAGMjRMLOtv4ocvUv078aLDMlMfOP0T9S7JKZ6Rbx3yYkHwsKW5dkd7d/egp+pLiT90DdxwduMp4ETL9+W1ghBadzINPG16krjIk0MZzKif9BOiVeMliFPVmy4qYrDTeqNuGbb0mdI85THE8u2OnRaUhuk6nDiSSFKgOKup6cGWqgaf4hayAH5RNLPqq8Uggtsv6a5q+PcMlqIMVwkeaHyf6xDy9c/MHlFA9jsomthDZESEKE4CALvMNokgYXCAUcCK+7cPzHPffS4kvGv9ZoIAQw/unMs3BEUyg1lpLoJgR2ECKFlIEYCcc3YSoYTjeDeFvBFVdKYyk3gv/YzG0d5MYcLokkwunFzl5E+Oc2hHq0i67rQorpn+9YyfHDyuw65b6OspsLKA/XA6tAvfSaEKRTyvshO2eaaakkVuJgTyG2iuIB01R+wHSgNGiKJpoCEboxVrA2jNHSW1tiUMI1kPwnyZYYA4zGHm/65xGQkFoPDjsIC4slsuyAI7roPvwnWJf8eUknSBAjDD5bxUoSm3CcSMiWJsOxIZw5BxqupUxOmy0cLAfKx7VeSPnkD98MQuggYehZgZpB0qxNoTWNQ0gYYVYw7aCDlFsnExv+wfeffPIRwZUViFVopesKFXXWtErCZdloTLa2x1M6hAoXpGySC9WBOn7Qjn8sbj6sJcKYHbWwF3FVKCtWqPsRJB2BDgmnjwdM6JE1IEyr2kELQ6inuiI4JSAAIfkEBQoA/wAsAAAAAPQBGQFACP8A/wkcSLCgwYMIE9pbE+eftYT/1mQ7aA8iAIMNL/3TKBCPwIcHe0AcSRLig3940iBE8M9Dy5IwY47s8I9ITZk478kEoEbgsoIvIMIbWRGnUaNCGgxUKpApwgkCB8ipM82gkn8llvwD8m/Zl6Ngw4odSxAqS7IEAf3zdlBnWBUJPQoMIGCgtIFrVH5Fy5cgp4EuwBYY+EEmKlQIEd8EmwNigH+A4MiUO9DKyA1H1wicpsNoZ4KeSnYpNdKpU4hnEwYtyFamTckFJQjUapA06YKnSe4SyKIvRAYDgSMs2tX3wFQC6x6VTTKacRgE7/ClENOpZoElBv+jSZDGv28jFYf/TXTGFw0lgc7866FCxRQLO6Yo21FOWTVM5XbsUGEhUP9/z+SCACcKHPRYTFCNRUtBbxjn4EHXxXRdhBBJ8U9uAgEB10h6OGjKg2hxMxBxMGkGyIEEURgdWHeB+KB4RyXioAKrDJFLDuUMVI2OXijjxT8/GhUkQTuW9ECO/4zwDwu5bPcgdGW4CJZm9fwjCEIESAlWYARZqFlRGGhJ1l9HqYITICoeBJ5A10lTh5hwlgRjigO59Y8dBh1iFHOoKMBFLP+chFA5xxiEyT85FvPYj14gCdExyvwE6U//KENQoQZRWtBPSKrgBzQuuEAmQpqleVCUvjkQJ5yPEKSMhqsS/8SBcXL0ZepYEZJ4kJ4QZVmQSrGSVWBBdhJUQp4jfaWkGo4GCpEyOU5STqOIYqpMoRdlK9BFmARpKVnTCnTStwZlSwgXLizC117/wBYsX3u8G2doviEWSijyFkSXQGpFhFZqIzXCZkzcyUiWMDIVe5QAu8SyIUFTVErQSScBaokhjmoK0U8cg9Xsxoj+g8nIh15EkAB43CDQKTih+o8Fvw3EARcF7ZCvmL8gxCVJGJKFmUA+DHQASWegeHOJ8jaEE3f59mxQCwJJZocvIpX07Um58JLkQJZCe/VBjlbzbTk5li0xuQntEIuSEjsasUDKCAp3pUEWiUkU38EJMEyv8P8VwdGZhVXJQBuwAXhBlAmksIvaHe54QTAYbBxcfIRs6QNfD/R2OSqMANfb/0wxRSx88AJoyKELxPZAhhBkSCAQC4RG6wIFc5CljmL6jy8yPaGlBo8HL7yDt5JkNFpzQHTC8MYlwsvq/zz8cElcyT2xQDlWsQ0wSRpCRe3BoPF9FcAMUcVAjkwxQuu0/zP+P+dTIck/twwBzPkjKVJ7hvuP4Gg5U8jPCIwRiECggBzPeEYgyBED5pGEE+qSmQN9AzOIYGZO+WqQmIonFqZNkCTXgYN6CpKgWfAiF2pQg/oI0pgR9OQfamjMQZQ0ggAKpAn/CEEfJCGJFAzBCDy8xS3/CBICKgQjfFUQHxWA8b0hDIGHBRHiP+bnvibOb4gF6cMocsa976UAfgR54RRm4D5KDCQYTfiFZsBDIcv8w2Uk+dCHDDI940TwH7PqS9C05LSB+OqDv1gNDGgzkMSNxQuFmsQ/WEGQPl7gH24I1vFiIoNYMWAfJzTGP/iAhmC0j37/MIb64re21AkEdAIZQwxWYBRd8EAXB8ETLAcSAzyFAwwxMcMV6NeEPwyBIAQcQRCCQAUDZMAAVEBDEAxxvircYgEX8heFXgiTO35weBy8ZkLg2Bc1OMIojUuIA27zlLAoJywj4F1ChmKUStDMFMBJ0D+UAIcxxKInEeuEJVJA/4KEGGJZORjBM6CJEx4IBBcxQaguWDHLgeACoSP5BQW4N5Ag/CMIwNhGFjKQAmRSYQYjEGipqgSTQ4mpSioq3qzm6Jt2bBAn59SmltwlEOcYpJJH20sRtCkcOKAgFi00hCUMYACEGOCXA6EiOMbgjgXYAaIxYaRApLpIPBFkE0fBBQ9iYANxAAMYGcjCFwVC0e/9wwDDXGYBjaGEbB6kX30Z2h7HAgk2XadngwOcW4cnCojgdCQkLQjN0DLCkQyLIKqSKUJMwBfgSCYWLAhp1gxgibOOpaFiwSxYGggTtHoWo62o4Qh6oMZimUlKLj1ck0pCVd/0sSSTBNE4BELOo/+V4a/G8UAzCpLHfwjnICBQrEFW+g+WIicKfCiBCviwT0rMYAZFHUh0/0HRhFg0JjywKkJYAVUpAeOznw2G+tTAgmcY9DqpoBeIUluQnTloTZCD09BwAjXhAS8hTHgkSe7xA4H8lixVmYi86sqC3iDKZP8IymrQct+wxIskFlBBLiq3tX+Q8R9jPest+gvRqgjkHQWhBywGYQYnrOq6F6VuSYpK1BYb4LtoDakaPGeMv/1jccJdlYVgQoz5kuUarYkVPLoAE/1CpGq+0e5REgsTloHoOoIiZEEaPBANhGIBGELosd744IOM6gX96QEfWFCCkLaioxn+hzhW4A+YwOL/H/39xxhCYBT9kaRDZChIdVfs4j4HYQQzsIILYyGE67BCkwTp8mmXTBD2QshxNYgmfEnStxwHa1QCwXRJuoyTY2hhIIydEpw+nRDgteMA49CAB07QgFbbCTlb/gcTBjIqF3xoAJ4AQRRUYIxcPGEEZTbG9wxQiF0OhJVoycQ/RtFAHOaLqGg2QLSHQFQ+gDSkxqjrjRPCAso0wB+EIMnyCJKA6iyFeS7A11Fs9rhjaCwsZhQI3sCygzfAp4IGmfUX3mDSchpnN/8AwSWQw6uD+OEfE/DgP7wDkUl44d1CE8ipNXAAHECi1f6gQC4mzAutybogo+KEKdiAaxDEQmsz/+DCNoTAWYM4g5YEMShOkH0UG+PE5gihdkeHkIKeU9sA1h4BC4wxhmj6iyCVoEQuYoECVjRgDQ2IQJZawIUTejzH6ThA0IbmY0uDZRlcgdO36iuQDvDCJjipo0FYGpNQH+WRF6hE3JUbHIEc/CCSUVqQhoSQoGng7xZvtTPIoLULdEIgreADoFqQCyLMjAEMYAMHOMGFfVCCD3zIBT9s8A8kxOTlJOnuSHAelmYkQQox0LZMfNhz1qcgGM/lwzM422o4KOEJlch97n0diDBQYG1ldqEL1dAKqHkim1RGiGkO4t6wOPqDCI6p1w9iuJLEGyKnM3BfEsRugViABZSAe/8l9lAJGPTgDhPggOShAQ0u+MEPbsBDIxoBCLgimO8GcUBfRSGKYeAABXgAAm/wBuIwB0fwD2IgEIYQDInXCm+EFf/QApYQCzOQeJiXAhmwS38wEARFUEaBDVAFVTIHEZwVA9AEei2XEDT3D+EgExkwEByVATKYAvtgRP+QC1XwC3AgBBhAAJ1QOc9VAjNgba0wA0JIgSAVDFSwD8ywN0pDEn4gd2dwV46DbwLxM/+ACphxWNM3EMxxTY/kOzEBTwUnFtVQJFYoEOJXAj3QA34wcmzABtqgDR1nCZbQCQ54LJmXCypQDpNQDV7gBQLgDXiAAwowBwqQAAngAIzoAF3/QAQWgAn3th8jwAyrsArI0AZigAxHcATbsA2GQIHWNgOdsA8DcYADAQGH0wfd8Ad/YAQFoT9jYAOf8A9G8Am28HLOgFUx4YEjsVEbJQ+8YAgzkDXO1YB80IC5sA9hlQGFkAUaVQiroA3FBREO8Hf4oAE+QHE+8ApReAHG4AtNQACBAHBHgQdpOBDaJxZYSBBd5yLSByfWFBaGwwZsRxKrJRBiOBKcUH29ZRBEdhDyJBaOF4eFI4erwA+gsAqq+A/bgGGvd21TkEIuZAUzlkIzBmh88ARPQAmUwAsfGZK84DyWAJIt4JGdkAuUsA/yUAgv+A9ZkBAPyRcj+A9Q1SoF/9Fm2PAP7/AIK4BLtmgEYDAG2PAI/oBQj/ANm2AG3cADOOkgGyUQDykP/3AEHNUJaIAGX3QE8uCJnSgGR4AMYgAKoaANccgAHOAHUQAA1QAAbhkInPAKryAKXRAP6ZAOdOiArdAKtlOSFxYxaocQ6VgSc5V8l4EW3Rcs0EEWMXURbFEXGlQQ1XcU+SgTZYhYEBFODNJvJDF5k8cAlBcLOyAOoHCKqAgR0jYQXySD8iAPyIAMAqGKDWkQsAmbCVEIA4GbOAF6D4ILbWYQv/kPvwlVIIYTRWcQMambMcEP/8APGbAPL5YLVCCduQAMuWAJKpmSfGAIfOBJQUAJJdlz///wnDNIBVTADCeEnf9gM8EFOyShJ+4ZE1RGZJEJE8nzD3NFEokpJkxGEJqZEGeBA8YzEv+1NwMxmA/SnyCiaQOhQfz2BgAQC9qwCjM5nhmAVC9ZEDwXk1XZBqlIEh56EMqZY6IHIiOKECGaECk6mynqoSxalQKRBc94BFmwUUeQAsAAkipQbwQRXCVRnzFRWwSxnwQxj114pKnSVzERjwOxj2NRZlUDALvwRy8og+MpE/10NCcYE+4AEb5YEKNwOCE6m0aRpRBwphCADGkqlm0QlquwDwa2mAh2OOxCEFxgoEd6CH+EFmnQp2jBAqcjENIxFuX2JHfwHyQBpP+wmEn/0gN1Kipcoi7bgADigAOFUAg/5IxZcIBtkKIx0Qa2SRCnKRAnShBj8KUEwZskqKojwaoDQXoH4XlHEapk0U8QQAK4mqskcKu8mgfxIBO7oaggIhLmiKQ4safMcwe9MagwA4AjUSt9UQwC0QixhRbSYWBIZhARNAAUUAvXEAeAEAfo0AjFIABuaW8WAAKBAAK6hgOccIl5AArxSgf0Cgr2Cgq6CgFtOqoCcQRikAUJKBD5UBIVwBdbUBApiBNIcJwJYQZm+g/6GrFoCrG7WrG8qqu4ygj5aq8kQAAoQIAiIBbqRBCX+Q9YYBDFaqzyMgAJAVcOElMo8A+h4QnztmBj/6FuMlF/E8ERCcGwBhFu/8CkMpEl0loQLmsMcvCQa0oQWUoSCZiAl1psLbENToADZuAK4bACFNANo2AG/bAJWMWLYWFivkENV9CJ/1CqB6GmoHAF4vC2Q/C2b1sFBEC3VVAFhFAFxoBo/7AbcgCtAgG4OFGhCBFkMME7hpRgRjGy8oICKfsuN4Cs/wCuLgsiDGezA8G4MHEGhRUTMfsRgDAR3nAgeHAJj0sSPDsSLoEQnVsQkUAQjxEJAkMQHxAmhfEPKEADuksDpjtPWBAOCCMQUnAOArFb/6AHkQYRIqAO1OAKK4gT6/APxku8cHYOP9AMzSAM9JC8BDEIAkEN//+AAc/ABQxZCJ3IiZ0KqunbBhEbmxArm2ybB9sgCQqUHuqKAihwCb5wBr4CtP/wAUBbrQgRbvFpEIZ7Tau7Kq2buTARBsQzEIHlEAJxDZBxEOjwD8XwumRRBw48tDAxu4Z7wAXRwatSuSXxGQKBCAdxBhhgBpkgDBUgDElQA/SQBAgTDjVwDgVbsP9AvMg7YgKxAiuQBPRwDh3iG+dgvANBvCvgCv8gBALRGSc7EmbwDwK6EQRxCcWgEbxzBkpwBi+gHoU1siRMwhBxxWhhxldSEuArJVVcEkU7wmhxCXSMEGg8EFCsV2tgU2ihCWKxIA6iBGssEID8D7VAEMtzAuP/BiI5cxBPGMcC8QsY4AEi0A9tvA7BKxDEy8Mkwck9/MmefBDU+8mpOhCs2g2ugDBJ4ApCwHAIQR0GYcZGscgIUcgwAU3L0xnjBghmYsI3Qw5HwXCHLBDDLFNQLKsH4WEHEcF8kQqNjBO/oMKIsGNjAQ7/oAvAYhSqkA20sGiqkDPLEwEqLCVpgBzHwQ1poAu6YAOMUMVmwHndEGnKZhCZfFX/EL0D0SGczMNYhc8FccQFEcr0PBDrsMrdkMnz/A/jJgVC0BmaMM8HaxC+/A+n9cyEfDQUTBCdYSEofBRSYM5hEdHhuyqIoHoEYcsEESYQEZwEsVvUHDw09Q8mDRGw/9p5AlHTAoEcDcEKrCANrBDTJIEcIF0QM60la3DU3xAO7EAQf6AItiAQ/SAQ3JsQTtANAhG8/gwRmJzVfYEwXJ0E/wDWrpDKEQAJtGwhnvfS/zDUMUHBI8jWvqE0yAFLnFVXTgYWeQwR4LDIat0XTzgQtMwXeT0Q8EVSfOwcfBwsy2d0AwPUU/UPTwnZkL1XBsENqeDTIqJkYGEHkqHOZKE0sPSU8HXUUNcAzmAGG0hn/2AL4WAGQ3zVYZ3QU20QVj0QUCAQvSAQpEAK/8AI7HDQmRy9SZAErDQIKxC8mVzPAoHJVy3DruDaWd0NLZjb/9ALYOC11JAJrlADP8Ayp//wAyM4gqfwN8ghVSKy1jZpB5p9UFp1UDyACyxjULjQIos0EHeNFs7BSHgCB45NEHUVZ0p8FKdw38bhZAN+F3DwCMqME8YbAVIQ4O+yEALBFgIMyYpUEHuV0RP+GI8ByQaxYPN2OJiWwPkyLIqRCAoXEzIEuwYBBzhmEOz0DzIEBGEHOdqHLwViAoWKG//AzO8ipAax2FBYB7cCAyWAKjW+KoYpUwOZEBqMNBBhJwImEBeuOAaRrQexUyNB2STBqL7hAS7gATg7HATRCFo+EGiHdwhxCOKRPPdJECm+MIULB+AxaTs+FqEyEMmjAJVWEMpMIdnKTWtBEJG9Kn4sK///MFgjUhITXRr/4Bx1ahBulxCFjhCLpq0C8SEMGiecyeMF8dcl8eQYLhBpsMBiIcBwcuYHgUEQUjwyIiMlmxCsXhAGMzi5EFnKoEh+CCRjceHVUOWoMxA9AD0C8YVHymSN+A9tDCezJhIggROTFji5MZlkoaBk0XwqWxCJne0QcQHcEecQ4aQCsQp+wALLgCQQlxBesCN+WCRjcS0jse4DMQK5kAgFEOuAYwE7VUEuoKCqYu0fFCELrgVwMQH/daSbThLfNBDecOmMXhLR/g9uQhIHPxIo3S5Hg8ZvjhAvThYsgDYFESky8TEk8S2Qcjvp7ixo4wX9ZjIW4AdsgO0x/+HlvrEKtPU4b6C5BBHjY24QSd7kq8IGP9OOYEH0YHHBTYETmnHeyVHBR4cWOBcHz04QmmWZJbHiA7PgoDYSr/a56wgTFvAEfcg1BPFuJ+EFEsYCirQMJs/rIoMolBIpmAApuqM7ZE8QSOKWsCutGewQ0hoAAcD3/3AggF/4WIAAi7AIsDwSgV0S4pDoCAdcXQjwfaEUryUTsyAQXIKFXIcTeBo81gEWiCHzCQHq2c6yLFsQAGAMPYBKJVEFdqhCRxI8IG8Q6G4Qb3C7YlLx3B4Ws+4b13cUaIflfdHfMNFaAiAAgNDxUmL6RjHFccIUgUkTdwe0rEAOrc8/+hmoA/8x+wVhPar/D2z5AFNA/gCkOcFuECNAYafkKqzT/RIzEsJ6NA0mCnnQ+0fR0WOBGdAAEP8EDiRY0OBBhAkNwhG4RuFDiBElFqRV8NtEjBn/mdA4sFKuGXyqEKryDEMYgd+UGJxiEMjABwL5tITYUs3BEf8M/QP2r9zAciNiCQwkoGUnnQLRGMjQ6l/OgcEGGjAgqSBNnzAFKjuGaRfBRwUbFGTyr6xEDv/SRhRV8FXHRRLJTfTR0e5dvHkVshjIV+/fjPUAD1bo4J9hhA7/MRRYZmCLFixG3Px3U8XAyVAhsphh0FiVfyF4/qNCcGmhKwKb/As2ZUqwnQNBD1w6ZCD/mCtW0QykUtp2wVtkgLVOaiCFIeJa/tEcMWPEiGDQWaNgWG9NtH85CMqYyMAgiH8WDmoQOE6vKQbe//poRzgiIYQ6BnoT+NX94BICi/y7VOufYr0AEMiOhz7QK5GCvhBIsPswgmcgxDpSbyA/colFBcpmECeXHir7x0LN/tGCpmf+uUW0jHrJqA+BJHHRBjAEUiTGhNgRaIiejvittIHUeK0TS3hCYwhxIljjooEUWyOAgazIDyJOBooSo/byWqtBLLPUMqEeHPunBC//eaNBLzAqoACBtOtIji0NkqEEGNoUaAIECBqjihli6eyfbcbQiUeBYhPosn/81KWgQyN6/wQXHhKdyNFHdVmgCquU2o0nYDKgiqfSJGkCHIcEA7CBSOQ09VS7AMSSGFTDxPIlvUxwIMIusLxkIBQEOiMvjmoFbIKBVkIhFsqCoaIngkgp5B+qDBhIHKnUmAE0P1mUiBU5/RyjCduCEIgKpoYAlNkggkBuihECIRAjBd0jL6Fp7qukEoH20EhViQwzIY+CHAoL1btKaWswYDNawgqBpCHIoUYgAsLAwyIc6BSAK35oJRoIyWmEXHgxwFtvMcJlIGwFGhmwk0X+p4km/IwIXCrKDWKyKWLJtSGLD2KwTXsjaiYiVHJubEtR3hXaPcTMU+jKow8qpRSOJHoBIgJjif/luVwsoQoYcMk1oKcgQ1YI0oN4KHsgszMi264gPnabitaeMwacglJp2i6m7yaoLoXWKFmhNI4eRqGheB7UoGzuUnogCrgQKG+MBMBD74x++SeQoZrLek9nDbJNnH+sAp0gZCFydO1/yMb2b9TxAsbt19s2oJPn1BjBmJUaXLegKpvu2b3e/zngAI1aoPyfUgRKXqMx+WPSrlgueOKf6e+TGK8lljt+IC9/VwuhXb7AvPCnZqAqhX/QN0CcJlj5V6/VJqIHIT1WwMvZZvOnauYRrJjMDR0oxm5NwxeW+DCRsWwPMMtYRrsiUoo6CcQvGUlLXDKSC4E8aSDNcw8H2ND/NPCM5x/j0IDAPICEBiQwIQdUyBlQ8AILBIJjLChBc5DSOYGkIBxJIIgweDgYFEXEDIPRXxEN4JzaGYMGKvREQtDxn47IomloGsgFMKLCpgkAS8uQSBMfEoU2KYNybqgYedpxAA1owAMRSGED3FEFcTzDF2bZDoL+YcF/mIINA/AECFQwAl7w4WrBGEIhhFCxtEUkZXZxFvqYlQLjRBKSQ6AKH5A4A3J84x4CYUwV/3EBGOAhFWtYQwMiQICEDBARd8Fi0+Llnh0oUJZ66cAEOvAXMh6EXp/kJQxeIAGD2CciZdLiQHwlkAO0J404YGMDFmADDLaiE3zIBWRYwMKB/3CAA5zwIBcI8YFAGmIbAllARH4wkHNKpALuqUFebPObFMRzCPFMASVTEAznxOIZMfhHAju5h3lVYg9PQIEu2igEAsxkCg9QwxOMBxgVtlIgG9jAP1xQ0X9AIiMDm2VBivkPAVFuggKp3kM2wIkPSmSXd8klYXZgAb5Y8QKUuEAlZNADGHBBm/+Y0EMmsVEN4AASaWAFHChwhW3wAoMDccoMSjCDju1jFpyYBRuUyodWtAINo9NIBBASlnf4wyCJtEsMvGqQdwjkEc4gSBAjkgF6wnUIlohOnpSgyYO6gRK5SARkWPjUGtbQOTOwXS4mwCaDOC4i5TSIRIXmgomaKv+WIA0pYIAATEJZDLIK6QE2d5lZhEzpew+JWke4I9NK1BQGPejBAPTIAWhogwuW4AUvxBGIYjQit4CIhAC88IDflukfgBBIKP6RgGMiTxRcAAEeLPDSN4hjFatARhv40YYjbMMAVOBDMFqxD5A4dQbSdGQGxkkHwqxDRhkhhREO8olP/CO+d/GqV1GUhQwMJL/7zcAQsjAETUmFEnQdb4FbYeDxCnIGhuDFPlKQgQwgVbE488bNBoIPgUABjV3wQyUKEIXA/WNnR5vsnCxKEGjIqRpZAqZC8FixDhFkpULDxD9KXBAq9sAPHmRDj1exjW3wYxX82AcVDDGDGfjPduj/msIf+cAHXnCBDdpYhQLykIBXmOAVRMBENXaAiR2EuWZu4AIoSAABPonDEJ3IKlZ5Adf8/uWsE8GGQsTqD1xgoxvzla8t2IoNe/wgHPE1ghE+EQK22sUIv1FIITKAX7qiwRIO3sc+tpGBQmThCFmQh6Y13QYSaEMg3smdQADwAk44oAvjEFjRRFG0V/hhHx+ipjECMRDQ5oUSHYVICP/hwOMJ96PAJkhKJ7JSDMYYL8cs7UAQW5DKikkinFgEG/TICWynAxT/gACa/7EsRk8lCJYwBBpmEJ3nIDmrnQDSgCnBC0vEG94GaDAz/sEPZBxkWQY5gkQSrZB/awTP/3hE/1jEmtZ/LHIgI0trnRG+JXn0+x9ZOE7H5MEPjGOcDqvAdo/ZwABT+GEEAHgDACwAyBYE0pKDPTcVKm2JTqTg3Swo8a0VstmOQswgNt/S9ewSwVP5WiNTYgAbZqGXQwyGAQNwQ5ir8YYhpOMKV5B4FvDi7Ye0odEF2bfVD8LYnL3vL+vM0hHyjQwx/EPi/8i3GJBxBH4UxOr7fnTdtyGPfVAiBRicbCxv/BDwiEcjRoPSQF6Mpb9naXIFiSDQ8+L4f1DRIBwkyAW4w+ulecebBBmTgCSjglxQWb832u8/wj2QtR8E6wJBxuoxL5B/k/Vo+U6I1jXSBlJo3fbYxa4Yjv+w6Sz8d0OdGcHfKT/qgxxfIzjgPELqxIWevt5UgAgxYab3hMtL+y4JGMjyMvJRhExNI8r+x2VqbBAFrCLTtqn7P+IskDbYXiCMIEHWCVNOJBAk4AhJTTcEws8tATuXmQj5cw80g4AzO7Nug4DWW4VXeAV+6QuBUD6i+QcRkAjHGQDp0wuUKIhV0hvwELqEOAQw+otSwYgJywjyIwjI+4daIK5sAARACAAlEIcgoy5kQIZVQEAS6MEEFAjXuwtGaJM5U4ginAgkGIP8Q4hMSA2CgIAC5DaCqL/6Gwge9EEfNLMepL8efIV4eIVV4JcLVIjm0aLnUQg/IEM5Sa4NbMP/fyCfO1hBgGkYhCA/C9sS+ACEONBDGYyE3hKAN3iDQAiEZ3gGOLqCVaADUFDEgViFKfwHUoAIrxMIiatCgygnsFvCiuEhIdiEgxiFh4DCHITCBVzABETAVThFEkjERaQDMFwFDYyCXfgKYXJD+1g8hZADVDqeO5CT1nGPOToI8WsTAoCPgSiG4QKEbDjBWRTBAhmIj7oVnsuLJzoIM4wC+BAHHNiGUEBED7gCKpu6bUAqD8ABCtAEYaiACnCGc3CGdTyHgXCGZkiCJICFGqCGhFCvgcBHgqgBWCiIf/yHdjoI+xHIiKAGEdiG31O7tqPEgzi7HNTBPLitXXiDWUSB/yjISI2MghdAATyggTogCCIwiFupmGIKxgbhqsHAg7lww4eQqDiwhn+QSYHwD4GIg+HKSYKggcHYFS2Zo5I0CCwoCBTwBf8Iyvugw4Egrn8AO4PgSZ5EyRcIhDN4AQKggIGQgn84B2GogUEYCFcYiH74h7AMS4j4xxWgx3OAR3jMiIA7hwpoJ/uhBgpQAp4UiKHEAAIQhysQgTyYgzwQAUZYBUbottY7TAi4gsRczCtghCtYxb+kgwRAACW4FQwoCAwYyojwAIMYRix5ASx4tgbhR1SxsF2ZRowISVRhysU4CN6ySVQJSUGAiIpIHIHIBmtgyup7CKOETYGQD7vASf+cxIhSM4hauIRyAs4wsAH7EYau/IduUEeF0EeDWKe2/If904ifEYjtHIgKsJ8kWIHLzAizTAhkfIhb6cCQVE0XREnAkEG90Mw2Kc+C8A/3LAb/yB32xAukLIgbEIjx/IcT+AetjIjd5DUkEIL8OyS90cR/4Mlq/AdaGNCB4EkK1Qtd6KSEkIIPBAd0oIVsyIZfsAERAAMzMINuaKdMoEdhEIgWFQjqpM7p/Af1Ui+yi4gbJYgbvVEVrQDntJ8TuEuJWAF3+IdsqIiCUAWDkAIh1QgkVQgduFAKVVKBiFCXrFCCeNK7oFKCAM6mlAhISKevG4gFYKvsNIgCSpK7wI7/f0iFAaKbgjgFMc3KC+XSf3jRf2BQiSAubiCIXzSIKVUFphwggrAbQs0I7EjUNegkhsCORk0DaSAqOBgFJzADW1CE2wgHgUxL/4OIHMUIPTiIUI1RUT2IdQjPFdDHJPhRukSCIxSI/NOEgcBTgbBTimjTjDqIAs2Sa3gidACEaxiIE4CEAb1QOTHWgdCEH9IIK82IPs2ILSAIOFA4ghCrczqnCPgboXGIDNXQghArsnIUAoGE+vqHVzUInNRWiHAIJBmIR8AObDkUOLULVnjWQ02Ie2iARyClBlgBJ/gDtwoHG/gH+8mEfzBYhOChcEgGFREIUuiFZHCCbtiEdfBE/xe9WBj9hyQIBzMoSFo9iI/VWIkAg3xghH6ghkFwhUw4BX/gAa+Sglct0GcdiOEkmZL5G2y5V4GgmENJV1Ywm10N2rs4hVO4WWr1VLs4J0J1hl39C40SCEiABIVRmGl4BGk4WoN4WoLQSilo2lNxiAZIUzRVSoXYJIGwAC76qYK4FVzERTZ9iF4kiIsQ27twhH8Av44yLoK4JSwBv02iW4RQDoTInoHQ27IdCLOtGMSQGOB8n1ZyLAqpA3zBDji5UsvNiBNsLJw5CMA1CPqgyX+IBPogiFf6h2g40H8I1stFFQ10j/Ncyn8o3V4zCEewWwnKixH7h1zJDw0aiGgDDP/vQwgVyt1/aN1RS0NVMdsSkAHCFYjzg4iRJAiF0Yjg7Yha9J4sqRPvaMG8YE2ESFxTEwiyFdsiEDxr5I+BkAbFeATvlSXOLC7KUYDBQJh/2B2BYJJGgAPixQi7FVy9sAcoGogWGxsoegSUEM2IqJUuqF7NNQgGLZiHYIWViJODgFyEWImx6Nx/YMODEDuFqEVUWQQEiL6CAN2+Jd3IAal/8MwtoWBZQhDJ+4c74Mn9JQhUCJqDwGG+7QA7+gcEIQIiCKA1sINS0t1/YAEJQOJjlLYaAwBfiIMMdQhc2MX7mIN7adLbXd2IAF3ANd6BmAZraBdYaRrR+gsSFouCWLH/FNYIC+4IE369RTDc4tqseGmlNfCG/fgkvv2HW0o6gQDgPz0I7hsIvl0qH/6HSoiFHggzAfmpY1DjgaixalBbiKiGamgyFiiccdLiifC5jkiLM0aIkiIMFrYLbsoIUyCIipKiu5negUggshUaYiOIE5zlLfmCkPJWiKhh9xjkgrDiQ/4HCfgJLiqIchAugqgGZEZmg5iEFZvkfziGn0AIMfoHIBgpXuLkwzgaCfhdOfkZAB6Lk+FebZ6IMyxnl4xhjbDiUBiAWBAjZj4ISiYIZ9aIeM6KiNgBFiiARDiTMxkMV7kPDt7gNgTcyyBnvNDaUkZngTCo+6jmf0Bghs4I/wShF3VWiALAqH9YBT8IhEmICYGYZoXwgp8AgEnAhHuWE+H6CRXgAwTRaMDIPo3w44Lw5I34z9ejUPA1iFA+lQ14C/d4X4lQkJmdCA1uLFeWaZGcAGCJ3ofQUjfc6b9AmLLgBALACow4hq0IKZT+h5ROCIiGCJEWI5AGCi9YMQAAADLbgFSGLKFW04px4eSxaTfcnTzuiHbFC2v7h4qC6YIoBS++Obuw3X94orzWC0BwCABO34LIvuY1sYTYGWQcXbsoTozQggDwVoQmCKn+C74IkX8I64QQ6YIok2U45nKQZpLG50c2iGLWiLLeiuT7gG0wNvew32xyQ3uRQ7tQk/9UuQ89vQu/xguphs03fogAGM42ljxs7qgieInL0I6LkCj5xVeDsGWJAAC+yCzRNohpnoQSYIHU9m5nTmsB2AUBSG/19uaIkObXFgj3jmb59oJqRuafEpAeQIAyzggvcWGG3gMmkEOsRQh1/e3Nxgjbxgsc/os2fojhPGctmYY4aITM/YczPGotGWRgNojE7ey9Bbyr0R6sFgguKutyaAleGIFyiG3Z9u5jYHGEKIf3lu+DEBAB2QUmCYBi2PFI2PHEeaI4gOI0CJxUIAROqBNWaHCJwO2BSMGBAAHzneizxWbI4Vy4/osUOzG+EZ6MCGwFUnKIwDmJoEMMF4geBoz/UPBliLBg4/HyDTKGHviJmCBtMQrrHTAGQ1Azn1jxioHo7vbuPa8GTDhtgSimKEhDjZBpZxyInpbyiBhJMTcVFxCtSNeIA38I7cDF+wBzjJBVR++nh4DgggCBWBjx0V6OGQCGIAntrPjzU4FxY1aGB6hzwuCOs1CIRm8TpvnAT0+IhxoIaBhuhNjjXs8LCA/gNlzsgxD1f8AChkgDzCEUPwfriIht0jY1ZHyDBzDxgaB1iP6Jn6CJYAAJn6jmsgataU8IXtcSJ0eIxSn2pjGBusAwhTjzDYxlwHjbDRzoBsYISHiGXHsIUy8IMVoorSD4OW+JcgiKXGCBB8DqWHKN/4FoiUuhAmMwiJiYgXEZaa+GZlo4ahkI6ICv64N4Av+G96aBAw9H+VmankrIpRO40FQ47IOA9YMw939g8bLmuRNnDdgg+BH/iRHYjdk4FtQMFKSIJ7g5dYF4gBUbEyYvCPtV6iwhvPsocJY/nlrQ5e9rmgqX3bvhd4PIjyeohBJQA0IRiidYqotXiDGOiTFm9YOfAjUgFu0hiB1ojp0AjSEwBJo48RGIjVsLBEMwhNkgDWcBhiowlkuJDSpIgdL4A2dp+4KgjIIYE7shJYeAA84vc+dDiCh3D2rL7ayXCGFHlcTLytfrxebW4hCZBUrIDI14e4KYgWv/hx4AjVtICP80oAJJuIJ98wl0KXxBERQq6P2B2P3OAZTedxZMHQgyWPXliIVcSAFLaHtwbwkmc+YdGEQ/QVbyu3WJ0DmMiEAKyiNu2m+UH2WB+KANQIXTZzGCeOzSBxiOaLaFCWA48NKCAAguiVSo+KfG4L+EKljwSejw4T8tDkfMeDglWMI+/yT9o/IPjcchkppkbCLpViBDhqpArFIFmCSRJBPe+jckoaGPwAz8A/MwBE0bwP5hdEjFUKsp/4A43BEsl6FgRZ+N+bfG6r9vDpc85ArxK0RxDkFYAHvAoQawaiFyWPTP1Nq4cufSrRuXAIqHb+zy7fu17NciD6/6fbgMbD2s0yD/ynCYCEbhfwX+NU6oKjLmuA5MOPA72eGEhLx4jTg4IuHBWBP5qFAa8WuVZxhn/rvi858thzVp/mti8o8k4L6r7P5XPKEtSZKqGBgic+2Cf3Z+SaJCBVgGnmDVzDCEJiEaNJKe6frXICHhr2XoMvjHyeH7ue3+zY/M4Z/bzPr1n9/vf20XdpXw0Be7XJKQVpkp848XECU2VwGQ9TWAWuel9x9EA3rV31cOdNFZZu3N8g8lCbmmQkO7qTCCISUmJJFDxvzzCxL/uAPWNoWN8s8YVS0QQww8xLBjH2Ms4MRDeSTEyEO52ZIMI4WM9E8KRv1zmkNVDJFCBpaMEMgCccQA/w4Pa1yIoXx0cbgWA3D9gwWacco5p1+0/LNeQnj+sxedfr3QJ1gB/CNAZI0NCKhDs7DBzDYDDCHWaP9kwCM5xrDYERVFIfSPCs/8w0NCcETGyj+k4jIXqXytg1sIPTZhABpBJDRCKx79Y0AGKVz30FDgiMphA5EwhSixxe53prF2BShXBC/oqWdCtfjn2mFxdrZsstl+FRpoCU2gBBxKxKKGaTNMegtHEMmK5ZXGRBcXqF+d+s+8dJWHC6mpVrVWvOD4ukW6vN7qEJcZdDKCMfsiq61/981ZH8NxEZpQDxHHJQO0/+DRFzdf/cKURMssSJeECf3ZIZ0BRGKsCX5xm/8QFzAr8c8CbpD7jzFU8MQRCZIUksJQthKFWjDH9XmvX0bGMEbAsgZBxRBZ8MTT0wYYMsIUxkSQ0IMWgzXNwms5jOZ8EOsHIgX6NSLAxNmK4vV/JzsE4pyC/mP3P0WoMOw/0ujX8n8xP4TCuDkQFcRQEPF8RMD/aFRFIMEE4leqff74Dzg3clR1BkN49HkQoeuc6RQj9BCDeX1Z899ZPiSUln+E0Lmmf2FHfEhcpch1aF8TIFD7P7o0AkJcmMDNlNxwgyU4HDS4MUIOI+RiiXaJqztwQhjwsH15atWbrR2gxsDSP0ekoF1CQjsEDBWhXz3CCOR0f49djfxn9j+hYJX/mRAJ2TNXJeqiB774oB2uQxRg+tSZtzEQQ+3hy4DYNZg1CE95cxGMYCy4LYf8IhYVkR4vDGCJtVhvLvg61al0UbmErHA/uIhXQsqjihjo4g/p+4essIe9IBiAh6GbAdZ6MAY7aDBiAaTTAYsYmVLoLiFvU6J/4NFEKDLsgf+og6hiEQv45SKEidNODuEWgxp1DyL4+o8PewiMq5ErfqJ6SCow5DeIJHE/LmCDQzjwOzQ9sU+2A4v97sYwUfSRiv7pIwYSYsV/7LEwTMmgIfHjEGnUwhh8OE0wqLfGYACDF5naFWYq10IYwhAzRMRMD1Ppw2CUbgqxyMs/HhTH2s2R/y7xwYybwGKHOkSSL2l4SAC+0MthrsUBhczjPxyWSAehhm8OaZuchrEft7wnP/+w0wtiwQcrzCAIVZrBDEqYkKEMBX03rEt5whfDuLACX2Xki/rmokoD7MQSBysNwqIjSzTpQC1n0dZnSGTIDiSEoIY8ZkLO8BUJ/uONDmnk2ApDmF/CTQJxcSbcLvCPI/6DARFNyCVAEIVcUKQTnfgHOIdSpVuJ4xZIcMYCIuAMmC5gE5rYwhYokC4bpI03xApjGOWZEHoSdSc9LI0a4HcGXdCPmE5FVC0H+Q/YqYUJfMllXSr2FdpFbJb/AICxqPqPKUaGlxAJRFlUM5GKPMQABv+gQAW+8oNVqSUTNphLCGhTlxs45CbiRJ851+LWwRK1h0BMqgqM4Ys/PrWIZ8Gff1anrQQ4cS5PsNhiNmYXyiYERHSzWIIcYji1zMd1aRmGB4TAVbpY0yEvsEAgtDmRYPBkpTYRBwV+kJBzZAYo/hkgLGyCSsISNwjws0Jp3CAIwrDCU36xIl/9gjv0AGoPjaViE1tbmLb8gw3a5Ys3HAIAPqHpo0XMg2c91AUE6KAB51mtWjaQELf44QwoeK0FWFCJD3YHLOLIhD/q0oxoYCY3D8nEP2owJ+K69XyDBSJy1WAMGiwmIc4FCzr+0VSwhGEtsqDPPy2o1v+kZT4hpgv/YyECzWx1hqy4dIsp8DgX64IFEzuYS2UKg1WLrWkcB0iiBjTggRO4Ny56GlF3u+sm+0bBAhaIRSJYAMRYlCgFVbrJRsLxDySt5XtgARWXweJbuZziH5uIjG0dbAA1q9kAEIaeMX7RnxZCBB3wjUsUlEjjh9Rxqw+5c58fIlaHBAAcfFkxsaKLplsmhNF14Z3xbiyXgmjBEfsJbcTGMdWpHiDITiCye+3gjibYAXX/8ApYZPyPAURBpCpwQy7ACcRgDIFJdDI1RLrRlzMnBNdfIUFCGgeRNRP7fG2+JHJZ8AxWbPgrAbXKNBrAA9nVxQ98eYRD7sywbPjlxE0p4mGM/yfM/Wg0Tq2osVwM+g83yAUaalH1Q945J7A26Ctp+fFZOi3kCLh3DRTIBR94UYURxIJ3MEvIfTgRY1aDIBDTmwEnr5AQmcbgXTFwhkN87R9b06VGDnnEJjy+Fo1DpErGLjaxDRCMGSA3Fv1r6oUoccRXsqIBYItAT//Rglm0oAVveu4wD/QP4iVEvtddyzEguZ9cZMt4drGoFSKzSIjkeS2hoRCa7t0OfeMAEu79gTiY3opWUGIfrTgUqiVpioV74gWJoMQMeCHxf2Ac4w/xtW73Awn/4ALbmSm2ldcceAPwAYgzcFfqsKLRAFaiEnvgAwp04d4GSIEAXOBFLMqRg/9ctMDadfG2xVznOtA/pCxThyJD5bIMpTeWo3VpQSIQpdELOD4hVZ9LA85UjWc+BHAJ+WeQccDvBjgDB9Nl+j+Y0HPkd3QCHOAAJxjACS4cghexpoQ2wEJytWytLqDqPtwgUHIrkz/wKSj8CPgQhfL8zypKcIPjZV6JCzwBBGloQAQIYYzSkWsKaniCH6ibf7zX/jyE0SUZIhydAspFudmFo/ncWpDdRmEGu+2HpDlEfjnEBeQC7clAD0DG1BGBQwCCWtRbvUHEKwha8HldA2ADGWzDCEFEMDTEzukcF3ABAygKG7QAH7QCHwTDNoSZX4icrj0ENjjEmeUdZoAfRDz/QoAlxAqgWfmRHxoAUQnEwgI0wD302/vNHyXkQi4kQgtQQkOUAEUsAcsh1RNAYJpAhIvwxTL9QyIxIaIcoLYgWhE1oFxsAB5xgqN9hQRcllzc3lcgGZ2wwD/M3vxVggyowB1wwfNxAANMALfAwCU0wso4hP1Mwj9wolqkoBNpwDAMAw5cgjWcQACMQSGswjZ0SUJ0wrmBE0QEHObxQQ+2giHwQk/sC11EBx0aIVhIAUTg2i/22sTFRRLE1T+8Q2bkSq5siZVZAjjFQi6ggB18g3udwAe0AC+8YRnMQAmAIzhRBPyogSHMAhfIwVfAUlz4ASU8QXupxWI0gxLZ4QIu/0VCYFSywIUh0oXrRQxg7AVkzB4HVgIMvEAPOB8bMAA0aAMzMMMsPMEXREItAIJFWkMglQNEBBJETJEoDMALfIEFvMEOjAA/rMIq8AM/yIPBtAJGzMC5NYQlsEA4Fl4nFAxYvIu2KEJCfEJCgIFPJgQp/INPBqVf0GFgJcQQOCOXnE/h8QEX5IJqqAY4PSVMXmXhAVErWMI+pMA25AhERFU7zt8ZwMF5JEaF9QnpxcUB2iOxaBaasF5cvIwFjcxawMWOAQhdON1DlMwG0h4M9EAP+AEbsAEHaIO7/YP12aIl5IIx7IIvBAAAeAFlUiYABAAg+AIOKEACJIAJcIYDMP9RFxCABXwBCLyBBexAIIgDKEBAG7ymGIjBETDDPnRlFYJTOFICL7SipMiFTt4dw3zCUA7nPxDnXIBfMT7EpNxEBjRn5xBeMFDC+bXCVVJn4VlnJqXAPjTnUm7DKgjOV+wCDqAFPgSZBnSaCXRA40VBHFhFDOxCZJySQwgihtihAtxjPurjQ3yXXKSefvjnP1wgFVVCCaiABPgBBxQmG2jDd+4DM6SASY0jUqlBLLTCEwDRGwTALiBAKCgAZ3YmaL6CHFiAjaHmDlhA1jADHSADBCADMojBdwIcdYKTJXBJQmTBVyjJjjiE3YFFcmLGOxzhI+CCDQSlERhBNzghNhT/aU8qwhhgAzb4wzswY1/gaFxkQQZgaQZERcCR4Q/mgpWxJJZmAZlmQSFkAQSsAryBhSx0gSiUggaIgnlqQALoIiVwYxUQQiC8AdEVS6Cl2lyMXl0IaFxkEHnpx5/op0NYE39u10OwAV3GxT+iCbZ4i1+UWwDlGREkKBtsACdsAEoiAyggQ0rKgzgEQznOALmsKqueRoXq5j5sAzOMxiG8nSUkwmjUJjNkwD5YgiVQAiWYFC5awqSoRSFABB3o1Vz0KFgEaUJgGy48YRP+wyM8gjP8gZF+QggcYUJgwyNE4T8YATuEgzOcCpXGxW3YxbHiaCFkgDzwAhrwQSfsAz9k/8E2ZMERmCm+HsERyAOprgIz4FF79AAAAIAAFKwFcIKHlIIxGZMoDMMccAEl+GArzCsLXGAC+Ue5DdpUicBcdKp8rWlhEOpakNe4EQuj+oeM3UdefsXkMIznQcTu9UVbmMIGxBgzrMIcPEQbfIUIhQf8tBI+JRV3wCTZ5QKw8oIlKC3T6iYl/Opo5Ei/HoG6goJdbN9XnKtaPMIRvsO32oAN/UM3VAUzPiG0LqNDmKt/MCeOUu2N/oM8/MOZbqkhAAM/yOYRyCYyHEEbrIIC+KEfepQfREHBFm7CvkIepIM2ROV1XiUakJ2vxoJrBChdxJ5fGNBaAqoL8MUHxAXJ0v9FnxaRJ15XF7hYX8jlWiwCG5gCJyToEFTBFdDBKoifciaEyanFyblVrmznNsgDPxwBMvzDKrDoP7ToPyBDGwSvXByrIWEDLnDrs/qD33UrhihJQsStXMRt3BaCGGRBClDCUVCBdO7DP+QsYjKoNmgDOo4GsPrgDGTlCASDISztdn7v0n6hl3wuWPwhXwAf6yhg8nxFazVSZPRjZOghsQjGyT7EzM7FA70HAzAAF8TCG7xBLIDC7P4DPzBvQiwnwVxp3vaF8orBQ1hpb8ot3KLwlj3EbwpjQjArotTLqUCvtNLFFoBFPDgEB3+F20IECZdP+bjo765kK7Yi77qr78b/bQa0a+d08KRwiTz06q9iyYn2BQjorz/1HuWqBQK8B//axaH20h69zHhGTC48gUYx31x8cWEcwgLThQU8Wx6Fxo1VMAAEwjaAghggA44Wa2H0rFwAW0Ik71dgKV/8pgtR67TGhZf5Bca58JLoR/ACckL8MEQoLyErb/D2sKTIA5m66ycDQxdJUOjaxUjahabpBV3cR6PWRSmDhS72CQHECd6oRQTLxQ7cWGoSy2chiiT+AxdUYEIYDyYEwggkAkr6MZYlhBGARXPyBbC5Jn4ai7L+h/I6BCXz7D/07Gtuc/nwqzzka75mAS/swxPEggRIGknWxQAI83/swBsnRCNx/wEBa4tWHV3MnF5clIxDFMR+dEYv2wVYRUakAmIQDcEq+LHtxgUnFwvtxgUk/0c1w0028+xDF4b4id9rIq8YtEHe8msr8gEiRlI8A3M9T3OcOFRmwKdchDFftExAr4Un4CFlJMSIZUYJlMASjDRfJgQyFMJSqsUyx4UgJ8RF68eO/kONeBwi/6LHzgXWOsSP4icEkEBVtwEEuCaLIsMVgMIrzMEApN1X9VLM/M5J3yNByfFD3EAZ94W8PYTnxSyOqQZ9ovRXnGzJ+PM/dO4/bG5ChAI0eCxQZ0HU3GjctgE/gEVRF3VkNDRYiNw/TLX2RUBUcx8M10WN7Atkq0VF6/8HCVg1aFf1Z1d1ViOD9f7DaZ9aQuwFWGlWScuJjMgFhYCnXTsEAcwyRKjjnLh0XeTYWEAE1lnMHejHcP8DPzfaWghKMZwBAXzlESwx8JJqmoo2aI928R51ZPRCE2Q2oEi2XSgjRPAiXXR28f6aYlM3dX/2Z6/CKyQADrAEX39FxbB0X8CJX1SqnHBWbSMKfYNFxdyBMJdFfzuEXP+DOk5XZFnQAGCdHBBCRQLCNcQBOjRCABzsG0jPV6IkKETzXDx0z/JrQuzwQzi2tmzNZasFIjsEEoj3ZjuExHUzN5c3aQObVRevet84jqs3e1+BB6A2Zek3hrwBWA34au93Y3H/ZF8YCERoVl4YQ3GDBZEzzD3/Aw2wI6IMACF4g0UCQhxYg0VKJgBggkiSBR4IAAgQgDg8ChdsAyPQAR0A2yoIcvDywzUXxgKId7Fo2VxER3QIwZ3XxYq6KItidVYXelaHNqKnNwmsQh64+RWQT0Lsggh2plxYFO8lRC3ndkKIIF24wFOvBaFEuUPoNhQh4pNjBlgGd7H0t9A9RA8QosVIVkKY5kOowAugAArQQGRcGFi0dULcQJYnBJfHgUXuwg28h0omRGKj5CpYrVpgd2IfLxBDxLGGcyEcwbGSwI7wGkSAd7EsUzi4QkL0gwjkwdw5BMflqFEXrxAPb4vO7qJ//zYogAIdYPA2cIE44EC+q6NYyIFYsPTGRPl9qkXGeo0vrAWnG9JN94lKy4mGghRYKJS29FNCeHk2ZKIhlUeGhScKaIkI0Dso5EGcj3Zot6iLXgFX9zgO3AAGdAMSVEAzSIEzVMDM81YF6EESQESL10VwyUVwKVhCAH1CBFfPJ8Qg9MMVXDsJkzAnk3jwrsIRPMMu7MIb4MEu4AGfCuYdeIInRIEnOAQKmNUNEIGi/YPEO4Suz0UAZ4agTMzBW5h/iAWGCMoufP3RtScJgkV6hA1c+smg/MPBp/1axPfLwuE/WDkgSFars7SVywVLX8LV10U989I1yAWidVhCdC4FEP9AIEBmZAK+L1xCHVCAgikjPfYoxtGjQwyCQ4RZCISDGfzDp38FuM4FPdDDOehBM5zDOeR8FNY+RLA+NeTBBhfC3vLr3g6yNy8/Nvv0P2CwOHS+SAVCFFT/GbQdCkA+c1NbeEK8XUzO2tuFQu1CpisP9wOK3IS/nFjkQ7RnWs7FgdjJV0hLpGPIGUzOzPi6WsQhRAAEoH//rA38d8mgwYIJCSV0OLCWwTMPKbqiGIdixoyB/tE40XGgr0AgMFBIMlCKQWcVKtRYkZFazEGDNCaElfDkwx//dmb8ca6CsCQrXhqk5krJroEEcKxalQcZsiNR27SBYNUqBK1br5DQioz/ETISJPKs2lbl2S5fvpTWfNjEbUIQcenWtXsXb964UfT2xYtRYEGBAv/pStgoUqR/AfxqnNjYYKOHCCMORBS3MmSNijN+rHnZ4CUdKEafoeBK2D+WwooOXBHOlSt6eiokcdk64csVN4WdO6c5obOEelZQw6BkoI6BGAhRSIhjoBMnV66Y3TZkG47shbYVwoFjCA5xN9By/OerbmaK0IG3d/++cSAadev8qw/fri44Aw07LHY+oTEgEyIhiygKwy1V/snmn/8GKsYaVeKIIw2NBLHMQYPmgwyjga7J6EO6LrukFuWUUwKLGzJRjTY96AmnhnV++y0jGvWoqZm4aMwx/6FmUhqoAh7/kSKJQYjaYqD57nPrBodqiQg99BJCzryaEKyrSfyQw++9WnypTMp/KiNnICy4dEicf5Q70y9pDAKkEVpAG8gzNo/7RwlN3KLlogrr4jMbPuccCAU23UplID6TS0gQGwbJhCYg/5kRLxodEi4vITWCsYJMnGPUIQP/yXKgOjb0i0z78JtPMvxENZSiWvhUL0ODkOzLxLs+DDGuH2EFDokBnWxvy4cUdWjQvvwcaNlENVIwURp+oYCdgVzJJBNhNllnIG77quDbu9YhqgLa/tlCUSGKdevKmk79NaE6/wmRMM3gcg43vda9S5Va21vzLnk1IhAJAvNa4/+fadpDRGC7FI0g2cYmbDauYBNlcCAGVfnFoIZBvZAuO/bTCJKBSo4jFV10AYcMRsxQxIx8cxootb68/efm97h9SZgbXUvIYIsTwoAiaB1SRUGOOa5rAcguWxqdDg0KcU0p1vTYLaJDaEwIou3CWCEu+TR6uYRutewhg/Gq5x+EGzDobYT9wiiVGOxqOiEF5SVQbb/SGBkvBeu9axPNdPFTF5RZYQWOFdgxo8AaDFpx5oxyfijnwhO6XFJuPb/LpZu5jc1Xg4Q+W6OF/kGnpmPZVJR11g3iBiU6DYoY3nMbG7yvpe+iJ3cuWSksZYMoJjkvHhz6kPa8UomArpJNzyv/GrfgWKP6f+C4PgZFnBjoD4cgH8i2h07K3C5hOKdZI83pUj8JoRKqwQxXVoA+IbwJTC01g9Ehuy6025hBIAHA9NlFQXbLSH80oidh8C14BkHUvCJokJr9QwhCwAUrcEER6Q0EfxW0i8Lq0h/lpQRTCTnFP5Q3kBUOhG7/oJ0dBkLDgTzCIfdglvGGl5EeGiSEdPFT9tzyjTWsIQZOUMQ/bDGQJoavH605yYom5xpG/OOK/wBDODZRuAu6ZSjZMshJvniXMpLPNSuon/1+cDyHSMFitOPVXVr4jw/+w24GdIjQNDLBf3SIgQ5hBQ9+aKiemMw9L6wJESHDx4Gs4Rs3/zwFDv9xClycApOUTIjcuIQwhOnwbQ5Zgw3/0UFBOkQarCBlXUyZEP0kpHr72U8oKULJaHRwgrrwY0YiUDJ/sNAgbpKaW6ZxxAY4wwxg2JoT//EHMyyTijUZyj9WYINk5OMhyWAHGGxgi8J9E2f/4F8NXEENyZ3RIevQ3PrOmARF5OOKyUhGP+znimb8gAc8uKNOhocyH/5jlQZ5ofJ+OZDh9XBxCQkiZDjYweG5kSI5SommaqI8RQp0oX2JoQtVyI3+TOMbcGglRy/qFoqK0C20NMgk4vICugggIXjoCyfh84BloBQyphhIB/5BhDO1Ci9A0IIjDOKFmigAp8C6y/8AJvAPBhhkAEog4T/eNtWEEDWpWbULqd5DS6DaBQBgTcgc7SIBEd40I3pCACe0ShEXDKCtFFGGFgYCBLdswC4qRakDEmKCRdFFOX54SFQBlxAY/KME/8hBXBnrFrjehaV14R1djmGXyiakIN74R71UV5NcxXWtWg1FQkb7j8f+g6eNgek3JMOYxbRKr25ZLEWW0Nj2lK4mP0KAQ6JqVYMcNiEq2Kxedmlb49YEoqK0Sw9dapCwJgQhFCnsP77a2HYtooLCdcFAkMom4QLOtXqB6VX/8YAp/KO2GUlASg1C03fVRRrWUA9dujCQ+tYXL3LAC3AT8lzI+PcfMjCIX+3/slu3tMUgFzguY4FgAWUU4bJuSYMnZbhgLhXgH24QE13w+o9QoMIgIN6pe6b7j0hU1y36zQhdE8KCEOtFbvMxa2NSW5Mu4FcvfTNIUymCC9y1Fy8ltiuLbfwQRmpEdhb2C4odwuS4qKC5MR0IHlw73gkr2a19ecJAMIzhDGcEpsowSIcN0l2D+FQzwv2HG0tckwB84SFamG1CNJwQM1MktgOJrl0QpuK73Pgf982Lfg1sEP3muYJ35utA4PGQ/XDBLehQigUogt1fFZoi4T0TgNsj07bBJ73/mPGZRHwXLxvkAw6Bg2YpQmZUKKDU0NBIjf8R5Uc+xK41OeKt4zJn/xGGesEMOC2P8TJZyFRChJZ+MX4wDWTnJrVQCbGrmAdCaYfItLNY9ou/HJJq0NSjzQ8xszn+Ueq4rAEOaQBHKmgQiDsYZAYjCIRSVMARFahgBBYIBGl+8Qs+reIfc8gIJugCbG0Dx2CFbrZdjJ0RWj87qcQ2CBtkrRkEDOCpT134DmElgPE2xhMDgbNMP44fg9vaPduti1m9fOp/fNsuAs9IqgeSiH8kghL/yIUxAjGSN1SjGpNYxiQiW1SDVGOlkwAAADCxA3y74RBceKpD4GwQXxs2I3euC8oPDhnC0FQjNK8Jsu8ysqkDB8QaiCui65IGzvyj5Kj0bvCUgdaalP/WLy6/C14VIHOHbPwfBYiFCpQxCS94AekDQTqnK2vUxv/j8Zcl+kCKvoMRsKAHgVAzvMBucC4tujEcSMiPHyIDIMQ9I49tEhHfhodc+4Voyu46ZMiaEbA7OyFuuotLv+BprSomwv9gNV3MDTe3HAI+PK7ElmMxhXIU3SFGlT5lDRL8SSSeIjuQQCwQS2fiK5nAAwE9XfZl6PdmhAl1kf1ACsugItwlAlNtACPZOnv73/8fXwj+3SOoco0kohJYYAoM7x8IbiDszu7u4vESYv8eohz+4QGFiw/SC/ncovjiAsG671fG71fSLyGGzz3OriZC6Ru8Bv+4ZJgi6PYWLBT/6i+r/K7cVoEL3AAIjIoBIS/6jK4B6aIabLAcvGAZbFAjWAoIWCAXAq8ANAzD1q8xEqs9qs7//sGvTIADT3AgRg27PIBN+MAK6SIFu1DbeIqn0KwvQiEUxKEHDu8fEhBWjkH6gvAB/0EIKeIBbFAFnsDm/kHs7o8K/+EVrNBogOD9BuK0HqJ5wFDbBMwurA0R2cshaowM60IBuisUiEAFvCAOa2IOFU8O/wH7fsXukO4OkY0BdIqx9tAhwm8KG/EhJM49EGIuWBE+CgnGEqLhBoLtREjrKGIF88IK/oEN/kEBoMEP0vABOvEhKuumhg7pIiyskG4THyIIE+IHNWIT/4HQIOxOCC3ADbgAr5jQLnyhB3In/PzQCitjEOnCt/DDFNXOPdgK8ChiB/EPBPNCEbnkAg0lvUSPA9xAGcQsGo/OIJ4v6CIjAAwPG2siEwdiISHw6IQwICkirFjAG4OxL86vPdLRIKpQFnHKFDbgIzdAxNwxIUThLkxRvPJC0/AikDRCBHPHDVCxgsINL3Jgy+RABRqyqG5KJyEwIt2wJuDQB9eQItBqDjfxGIUQrTAhFzigw6LQLpwQVjjyVxRxy6irMWjg/V7v4eDFIlESOKCSLrAKq4Dj7Wqih2BAJv/BrmRvLbVn9vJxC1thCiKyLrDvAZHuEymPE58vIexSGv+z0ejY0CCiANIGwgUbIxZhCg7Y5i4YMasUzCBGTVlQ4PUGwhUTIjE7UiPGiyb74hbvQsVgIORyj7F68R/IzS6qzqzILiH0ziHUALFi4RjLq7wIMyGCTvqEbhKU0ROPIeiC7geHkyiRDgHpAgF70yEP0C1UgAg2szEgkyIOMzNtSzINIhYNwjE5My9Q70w+U6uczFA0Mi/Ygy5cE/nyUCNUgA9YIBMfsDaLEgKVISd7kBPlEABgyuMCQAD40+MEAC8DEy+WkSj/AfocogiI4CX7Ygk2b8+gavauMzTapD1SBTIKUTPEkjtrQvfe4y0Noh7/wfcyQuZ2USMoMyMiKSH/MKEEWOABqO0vqTEhWIoPzosNg7AZlW4SCG7petQnp9Eh2LAgd1A/HWLpjHTpBAAEyNAE7aIMEqLq4NIhFnRFj+sqa/Hg1O4ABmIc8mK7PgynECZEYeULOS4vKtDicisjOlQveoAFdoAhH+IY6xAZy4EPKkEZAnIvkTHojPKm7FMwHfC59JMxAqAYGgEQJkRRJyRqWKdCEocwfGEAFgEcKcJ1/uFJXcwguM2paoI8N5Sx/K/i/OK08A7v7CIOUFOIfk8zurIvtPAf1qvj/mEEltMBaxNXR0DN6vIugnAe+4KlgnUgjrRIDSIAOKMR4gAQAOEMMNQuFDHUAGBMqbTa/0BVI3zKBSo1IXKxL4IRLA2CJOMCBA7TIE61Lp5LVe8vuf7PIGDTLxJAVrdOL9ztvOKwHMQMRh1CBYJhIKokIXAzIwC2LuLQC2yK2h7QqJah7pThGPIUE1jqssbLDeIxLp40IbjNWQdiF76A0rKTO7kuqVzAIsnsH3ygZO8CAUjWLogMy0otYylCPO3iQw2lTA3CD2htZHag+TIRRhvyGGWTCv5hBphThOLTLnoyIYiAAPTCYu1vn6z1ruKK09wjBdM1LnCg/ChiXbswtdblDXqgVh/ivG61Vg3AGKjRaPHiAZAWL/KVIh6wHNBq/0LuaSsWL8hVhPAW/9DULsgO2f84QEP9Qi7vwjs1o2bxAqlQwQUo1lpddSAUZhynwG3/YXITwhIMwflqUxnSNi44Vy8s721DFxndo2mPC9LObrfq9uB0rCYYcQ8cgq1UlkvjonCh9lfc9eB2oflsk20NQhlyIOf4lQ5xtTaPcyAua3MTAlePNi7KwXONFGTxYxZstwvx4WRRCjwJd7hQ6nAdrl3/gW+D51IfogMEq4YKBU411y3iMN5s83np8B8AQDEEoBodoifTdgS4sBOGdk7Xl3IpIrLeQHVxyh01wAFwjHrZRPQMouLUzmQzIny5JHvbqiESuC54IApGgGfpIhY64R/OS8zS9j0dQswMkBpHIAf/NjhOm9ch8vcu9vQu7jG/7CJcLdhQLHIgHth6H5giIvg9Jtg9ZNiG70ICXJOX6ioj3Pa8ZNMQHCI+PfcYnQ9tB2IEWoESxnYg1pZWsZhW0cAgglZGB6KJgUEjKhf3DIVaDcIkHQKB4WOkBuIqVWBEk6rOIAM622odz8RjuSQ0caocayK9EqEDOiASAyQvanNo3dZzM3Fo43QK1GAG9JeLDSIWduC8piBsm7iJG5kiqIAKUsAgynKSHYLgtvYKDcIDYaUU4EW4PG+IcSqPzwS4hBg4+jiCwi9e3WIJSuAC8hAEiiFqVgcuDeZ9M6IVwtYgjrEh7eqRxXYKuFBOH5AL/wNhB45xBJrYILy4E6YATg3ChdEgCFJgCAbyg8kZXwfCqABgF4DYYmn5Lsb3IVb5lemiABzXCmO5L2q3MbhKI7jVwiqDl3Ph3kYgFp5AHIhAHAhgAdCBHDYP15K5JqagNsf2AanNGLjQ+cphBKoYDapgILDYvJA5AAJgBDw4IahgCIYgGEYgGDpBeP+ho//BAP5BEsgYmcnZiT3xDX5levXWCh94jZXsdR1icOdZL3BHn/GPD9RANg2CqTO4VkeZIi4zbMshDoEginPBEMyDX/n1vPjAEGJaHKrAGMwrpL2ZI4Lhpf+hCoBBEtraiwciroPWreHiD95abPlgBLj4Af+ALhB8ARzQARx+YQFQYAxQoI7gA84+tT2+1agzInC5xJQfwpH82CBy+Wkvy5YPrgX+YXfzwq761yCcMD6V4QGNoa35lZPlugrQgAqAYZxv4RkkegqmoBWw+R+CQZPZOhjaeiCaQBLA+Iv/AaWRwSDAgAzAOIpjwRIs4aYHcq+rAQDe4A3mbd9a0i8GBQW+wKHbGDK0tTHM8/5kF16iLbgeW8kycCBaYPBks6nL+R9kU6ozggU09X//IRC4j0ziGpvRwL9fm6aXSBx2oBxs2xB2eyCC1qNhuxAkYZyHoLXjOsHremtu4R+a4A/ImIoNwRJ4IQj2Wmzd05LljSMEZCD/6kFuQi2VNaKpzi6NE6JLgYOtXvwughoyJhE+ZEq9lUx+0RteFu2P6aIFWoAX9vq9P/qDS+C5NYIFkHltAwEt+mAgPNogqqAKUsDBwWAgrgAYAmEKdFvCE6IKwFgS/mFrMBwYcJu4M6CZBkLKLdzCgWGjuTAIMiAIqmAGJJca1cAQ+OCYa/UZAgEctFNE86I6B2KPH8Id88AvTAG884KH4wph/GTHfdzSUzEu7NsheCEXlvghRmAGHFojQF2KafUZbqEPbqEKJMEQqKAKDEAS3trC/6Eb/kHVA4FfvTiuO5oKZloSbmHW/6EP4MLKiRsNyvzXl2kg3OEf3EHKNfwh//IcyQu8FSxBrZ9hIMhBF8Buz2qrdN2iUqWzPab3PRqthm28q7Asl/ViahvjV8+kANw5d6zgMjG9PSCt04+8qRuZrmpryByCD3Jhr6fgCIX9Fv5AEWIdLiiiiQDcrf9hnGnaFoLdICh+zGFbEprgFpR9IG7BHRaAB2Jg1QfCADJAuJXXhTuhE/zbGChgDKwWVtpBhCRTQi9dM2prxmqLsd19IJIaP2TgsKI0gvIs/KiyJjrbIfD2vOiK07t5IFZ7IMRMv5ugChbeIeIhIWzABgyiCazeISi+1ivewTH+14Xd7CnCGWLAHci4znkhIQqeilf+HywhtyUBA8Bh1+LGWP+FyiC+vSYeXSPkOXcUrOZFaDvBEBwCYQlqK7Gk0j2E0OcHoo6B4wXEPan8iq8cwAT+0C+QPhfUQAXG1hCq4BZCnVYPXCPIwRekHDhYfyBCgNn/YRTGwMTdwcJDwJoGAptqAgquQByGwMHLnLXN42wHAsINwBKeIVV3DebpAvAfQub/QQNEAC/I3SAc2+ZxigVyYOf9wi6b//5Q9Ey4wKdrdQaC1sJrlaBh+h/KkqjOCz1M3C/wZiDshgewG0kWIAbMIBkA4p/AgQIhCHQ28A8jgbckSRrY6d+OKSMEUsmw71+wGcGMPQs05te3f2sIPvinhaDKlQMXsXypchjMmSv/Z9G8iTOnzp08e/oc2EPgkp83Mf174IVgA6JMm+6U4BQnFzZchuQCRiUIFZY7RqD5h8ZQRYLlWAQiyOMnHKLxVvF7OU0gGUV9QrhrAgws2BFTvv67mIKKISpoCBuqgiFOyZICi52MCjmy5MmUK8MM+g+q5YHLerpxA9PB5qaaR6sUV8WduH8pePHK++zfs2CG/lEK8m8GwSkqRtD4x8qOQDtpKLPCOYSlk3+jYvDggXdgMNq4qRjIoHUgFWBN0K0VyNi0+PGRl5I/f/MRz2sEO/sEslK0SvMEBxAVwHSJBGsvu0RmYN9AQvQwxUDGyPMPOVhBFAQfagiU0gjkgIOL/y4EgWNahSzRARM44Izx1z+1DaRVChkYIJA4GfBSRTFrhRdeMegxxcWMNs6kwo0qrVHLP0P9UwZLxe0U3kCOHEUUfKX944B/k0USyT8BQEafZDVOIFCAAilhzIP/TDHYEQOlQJBgY6lR4Fk0HTeZHRbipAs4uujyzBBVbIWbRbyI8U8GGQTGlzGBLDZQlTDtYplMherEwWTtEDSOjpCJcl6QQf6TA0FD4iTNSrSgNJAX+OEEwz+gFcGSkzT58VOUktLEAEtKrCHEHQ+qMUJWlmQw0BAPCZTclwKNYAw5M+KyE4j/LFBFXipddKJFVAhGUSBpFUmTl6+uVKNklArkw/+j20J2AFGqzvTjpaO5xxOqBJkg30xYtvpPHAJxA4gqArFHlAkmCHSuTrmwxACr/+jQ5T+4TrvgP1eQ2Wtylgw01rg33aKdRddB/I9WQQRhCJojLDAQtq/CeFO3DMwblQaVJUDBq+X6FG/APklxHgwymGqBxT7TtEAPOeaWnUpt/IMMMAb4SsY/VVTxTyDF/szSL+IsqNV1wZKY1bQjqLFDFPb6LMoq41Xys8lUE9SFKDavzVO8//zrlKsDAfDFP+7BhwI3VA8Q6xlr6HBHpiPwYUkQKGYsUBb/bC2QL8be8otw/7wJ50CY64LsSp3npIubv5AjSdcmkuks11pZ4uD/FMb4UtJSaos387eUGfrT7E3pDndlWupUIE8ywOBuBy+Z4Ipkdgu0DHz/4NH7P4IvYExFI7TCS54wDeG45mk9x6ZOnX/++U+d8zCnHSBKkteff203rerTBsNXFIFY/k89OvG+k7j/uBy9zfAvMjOj2UBE8wqLbYokaWiEQEpAENCshG7oYVcABUKD6uHKEAYIAjC0948OhqhjK7EDK3CRFoLgwg7lM034/mEHO8TABn+QRCHyEr+tqEQr0wIZX0YQhU8JBHcXpJoLNqCSAhYxNAMpBU129hOb8EQLX1igQACBkwLoSBkBjBV4MjiDB3EwT6nLmA5VgjkU4kJD/0BW/wubgr+BvHA4EcDAAsZwQxCe0SIfw4pWgjEFighhIPojSKZs9J3KoG0ge6DdaI6BnlLIDTJS3EmOhmSyUdGEgktsygnuQBOWrcEXPQjjCDphgIkJRHtbsc5NhMM5gXwOcz0Z4Et0AQckgGGVNPFjVoIASN6IbYgEeUEnozI0mCDgJ/gYiO2OCRMnEoSW0FTJJKspEE6uhAYweMJAFqkSDkygDnCoRSnFmEoShvAfZVzJHnmAIcmM4h/JIwoJYGIAHebzY/wEmRpUoIbXrSUuAtEXZOY4GVMIBIlrU+Iz1XIj0VxTINSspgMcIM23dQubM4EiS7BUzjs46JQd7OAHU/+Zzw/SREyTicBwZvJGluSJlX9Z3C/76EM1qKEH91MJJJJpGQBCxgVN8WJUlEiZ5Y2nFBqQpo5AOZ5UVOYkneFiZCZKE6D+gwEKFec/4EBKB/2jFQbICxrQgJtcDAZF7SQRivaoks7hz4QsielMWFHRlyyOJSgqqeI+xheKjOAXKjFoU5RwOZ/YUiBE5SgxeWI3AKAnUjpiwUDUFZm3CaSSMIkGTDRZGWlilSAQ9KhKFDqQNFxCBXywQm4socpgVGda+YQJbkAIEwtZSDhx9Bx5PKi47QTXEjPgC64GJRD9SXUyeSOIyx4Vrn9oYzPf0IFAJDgaH/gEu44dD2adMtr/f7CMJp2yEQDDSxAmwAS1NmGPBZ4wghHMALYRUSeJ2rrO2q6TJrq9HBtVqAs25ZUyf/Urcb+mAhUYgwf0WW5kQICCmfhvM9Y1JkEsKx6hdpcmsSAvU/Tl0e/6JAFsUwkGBmLUjarEb5xhiVVD+48EEqWrDPjAPy7xD0L8I76wDcY/+HBbmqhSIHvFr/cSe0vgKBmGSP6Hg1XSMIIYeSB+NTAawoimWPxmIE92SoRX8lwbaTGAxlvbQ1cCAoJYYCxpfskyLzjeprhrbY16yRt6wIcRWKETlAgj4v7Bi4FMjAIUqEITqlDomP0jHP8ggEDaGgLJuGMmuMVJlQuMhq/p/3QEPd1wTp4ATmgmUlKU9cmoPe0TFcx5XOrdqkDevJIRxEI3fNBNbgjCVnKskKD20J9n39EMgazgBv/AwT8KIZBIEyWFO6n0TEpqHUxr+riEFUiXUb2SC2D7PPCCyQlwYkWBuKQn3lwJi3UEvZmsmiiZEIiGN6OCWDwhR0Oxwnw5xs4m/EA9K9GDHlZCj0yY4R9NUPZM/pCT1azm0U4pqQFKqrQrq8EKFOnBt60dhW2zRNvnKdc4tMtRujnRqS9ptUB61pjHEsSoMEHEQEqDxYGM7UYuFUgyJ2GZM+MEwwRZ5ptVLBAQxFsgrlXDn4mcok2oxB8/aUKyYaIIExMEA/9bwAAGXHEDY9NEe5W+dEklbgVc9cC6RNyM/0QB6w03s9TvZooDJVUKkg+EDwNhAscJkm6C1JlqmiWPoYwCmbOI+B+oXckXQPCCXNhaYYh7uEqa0Iyy+8TgBH/6Tmow8CkL2r59fbjnPy8WXKkhB7FArFO8SAScINWbp9a461niTZNPxg2yJ8gaGpCN199EAyD/B6VCcYKy/0ggdy/83lGAeBDEgg8ssF4rLLE4FK3GHaewxz/OkZMksMQWM6H8TfSwAktTefyKe3j5Pd8JU46+9HJ0SurJbXrLlFsn9NA9SyD5E57vZO/3IYlA8r4TfXdBpeYDw9BUwCc7BOFZQHL/KY1EeAOxd8ZkARYAAnimG/FlCIG2cAORCT/AExVAE9w3EN4nHp33eZ9HBerXGyBSEscxMDwhBwPxfiuBVATBBgLRepbhgPtzEzUIGaClSa5FHhhFEOu2f+P2aSuhSXkDgFHBfzPiPCvhBCT2DyIwEAqAA8FHRFDRgDWxCI0igRawAyygbUsQXxFRVgJBJuKgdCohDDDxDiwRdZKyV30VQif4eQ0ievH1G4VEE4tFEFo1YeRxAa3WSDsYGYOIE4C4EsFDFPgHGfM3Eyp2gzghif/3PKbBCXAzDo9SLhowDB6ghT/BBo2iBCAwgRbAAq2wY8VFCYGGdP/AhsJQf+HH/xJMJ0v8ZjH4hYd4aAnBsIdR4FKSh4kqUWY80XbjcYkQxBO8Uy4+uBKAMHM4AVqQAYkzoQDZpCN0BxOARxNfUA088YT/UF7ngQfnxiQCcQAfpwFN5QER0ADxqIA+ohKhJhAKNQAvgIoWMAW5wIpmmCuw+Dg3EQMCgQREgTE0oYtONhBbIH5SdodKg4fikErA+DWcVm1LxhJ4MDaM4QctIBDHyBJAJymsKBD6lxNxtIk/0Vz2lxMrSRQ78A9vYC49sYDbQlkH0I6i8I7xeHu48ANrMI0wsQg3OABngIoqwAKHMAPF1ZSqdE85cW03sRw7cQr/EIcrUZD/EE8q8St8hf+HKfB5vyh6LBAFzPYS2oYH7NEAa3AcfoAlv1MyBKFjnjZzhUce1QgTL7YZMrktO+CNLjkT66iT7egBiBCPDWA1VXAC6IAZAvFd42YKi5CPqBgIuUAJLFBcwZAXX0kZXRkVHqiVAzFwLPEQJyiWD5cCSsMLrSB6MxAFx8E7SwAC13B7a5AKFACXAmEwKiFE0VOJi0gQCsVQMPGJNxJnkJGNaWkjO0CTK9GbkMFya3EPlSFZL/Et4/CM42CYkJCY5CAOuSAOanJZl8IBLrGSHHCUqBgLuRAL8sULyHYQWxkZaMkTkyYQ07CQ/4CLKhEDV7kSi5OaBiCWBUqgBEqWXxP/C4FAHyNBEJWgbSwAAtxwew1wCo72D8bzkdGJTclIEHqJCoMJE6gSmDpyjTARojOBiKahXjT5BiU6GtUIBzrgBitqjAIxZjrhHtiiAeXSDjvpAakQj9jwDLnAB7nAC7lQEcyodwNhCqawnj3ACxfQlFfwEPQpEFhqGexAEFPJEtb3D8EGE1o6EM5ioGf6cMBgkbLmC/SxBl/2D410AZUAAyiQBj55oQPRArzQAn4glyzhif+gXeiVXdoFjSqBGdNFNUK4E8dwoj3RCjtoo5bhiDQBkjOhTeH0D3vnl8UUSpShAeLSjhoQpPHoDFDTCq3ABy1ACUyqEgzwhZM5AJ6g/3x9lgvIoGg1Nxr26RP28Aj7+RMHiqarST/xFQuwMxA3GaeVsAeVUAIgEAeJCQkE4AdcwAssoAKH8JHQlA470amu1xlG6BN3BxkotxJRyBQklqkzEZgtORAvKK6PCRPXqRL85h8u04ntWAo4IKQNcKoDk6p8QAkgyYzqFWiwygFPOgBRYAxJOgMZgQQXJx4/sFwR4KU4AaYIoasdMhC/MqwHWlYWyQLBgA62RxDNegG5AAMgcKfxGAHiwAt8MBFagKQ3Epw94TLh0nswcQjnkZwz4Vo5gK4X1AEcCjz/gAnPSTAT8LMssa460Ui5MKeRkRQs8S2FKQr8Go8VIA6HYP+SPzawuaB/DMAAHMABnMABXBALSRoLhiCf1hUBCIETZKoSDqoSvCoZdEsQBXkFuPaxQ9CaatCUzxBH34ACTzCnKFsJMsCy8XgCz2AMU4AmU+AINUsejVWcP6GIP2NjODF8x1QgfJmEn3oe2gahF3ABMmCuOvF2M5FAlPItTaW1/ioOE0OuuiGQE0C2HDALHMAA1voPy9cJyCAQOEMQG/sSohlXj/BGy4WlUoW3N4EEj0BQTZECBXq9BMoLITMDJWAMlnN70YACBZC4EJoLTACtEfAMsZBgOhVIlSuQO0GoMLEBG4CEPNF7m2sxMKpxeEkTiIhySgsTf0oU4vquc5r/uioAA7xQZwSMg3EzENyZtf3qDDZQIy84d4DGC9UqXgwwC5zAADdYa3zAB6tgA/8gsU1hVzDxHEzBb9Hwhj9xvTN8vcDgmk1JCBiSmHaAAh9QvgUgtUnKBxIQX18TdjrVCbBYvSyRjORqKMQoEDHoE4f6EjeLbRbkE7V3E4uwiTB5E5MqEQMBGk84AEYbGTwntajLvjAwAI1iVO/nDTCBcwIxxwQhGk3lbllLoQ3wDeEQCrDYCdzIik35irPABfvABVzguxdQa60wA7zyDxlJkC6lqw75D8w7EFk5ENFLE5BwCv7AA2Raf1jpFDScvUEQX1bwBCjgk23Zwyl7AYng/xqOLF9LMANWoGfThsEDpGFcgME+EW6jgUT+axr0ChlDu8Urwag7YcU4MTC/PBDGZGHj+A+mFRWAR4Y4isAyoMADsAhlOwsTYB9EAAMB0LoqUcc3Abs4YA3ckArZ4A5XsA0ZQAljlaoCUWszwAJ8gD28YMhG2sgzwAur8AeS/A96exOa/A64oB7a159ZOrcCwcnIUr3t5hOmfL0bIWvPEANrUKE04AYXsKew2JRNWcszYIa4MgLxi3c3MQGV8AQ0AMXjkrnkYcyoRs2VcamXGBUyaVl7AMtAzc134AdfaLYFMwAd4AYBYDdY5CpzXLUr0TYCIU04cAmXgAd4sAtD4P8W8gDJqVrStmZrrTnCHNEJQ9C38wTRCO0TmsCfB32x1sYDXRZPCP0ILERP/3DCOkEmKTAEfn29vHBlwTsGdnAPDYALgiAOldAKGNaUZRDWtTwCtswL2tC0afcSlZALrFxELkBUNW0Zq0av38oUyHwe93sTaKPF/UKFPSGTMMBx5CvUKkDUaMsJ2gANVJEIH4AHkdAI0iiN/yAAXpAUUa0S/yIasOsAOPAFb/AGILADubAK8vwWGUAFqjrIJ1nPiteUG0EJZAI5BzMQNUcyRKEebv0PyssSIGILioBwBLFLOPEJRrASyLsQwMIaj3M6fzLDPvYPllAFxpALYpsbJRD/1gde0iMQDJawD0PADAJhXf6XEwMAxF+2FEtsMeMF2ptx066X0yyRo5AhgDPxnB2mbVIr1BbQA35QihyA27zABbPgB29gzo1g440QCQFA3MQNEyInUQPQ3F/gnIHA1W9xBPwgBhnQCbXh36944M+XAUMAyTCxABFQ3jBRmk5BCirxB0ZACvP9D/TtEz+wlcgrEFN+5qdzvVRwOJSAwU1p4Pk8A5AN2cVlCLvCC0MgD5xgHxGeEweQAH6Qsi+QSIzYE/EgEPr7EgpFVI1lGlr1eqgNE9B8E6jFcv1BFDJwAVok2xcAA7TN4hzABmwADbA44LwQCzTu25Ew3DvuBZNg/840EIPL2QUyJklcAALNbQFvsAOYgQz80AZi0AZHcAQrksQHFtaWYCJnLhD3fbwCceVXvn2j8eViPhCkMIc/geZ9wiv7fb2GMGuWEMglXWuQXda1RgW88CdRvg3bkBEqEW4+4DI9ynuBPqdRMCQzvRLLNZQ0oV36K5M+7ZKmPS4CDMYzsQgKdek/MTT8OxDa9uk9IAelyAmkPgu8UM/1RcK5EAggAACTMAmvTtwC0Ai7IAcKoAAJkAD+clGlIAIfgAmAuQM7YAGYEAur4BbBLgbEngXyIA+8IF8mjT0qAcm98A9tqCNgwA6KsEufcO1O/w9bLhDYThPW7p83kRwmIv/ltjED2NNnjnzuTYk9JuInUo7WXoydTMVUo+oDc+AHuVAJGYcIGIACu8CEvrATadAjprHh4PIPpRYVNAk9HW4ZmD0ZaK8SgOdN2hbiM0HMx80TxxjzzOnpKiDxpViK0KANK4LxlFBrAvEgM2CkLFAO5SAqkUAD4qAAqDAHKQ8v8JIAA1DzMV8E/BjdoAABEIAMyHAEYrANR/CLM5DPfEAm2w4Txjsj2OAMlPcJkfYN3QAGYGALRgAG68BC6mEHnDwTfvISfuL9VLARvMA6/Cz8fNAJyu79WZABWcD+/LAK2yBeLxErGNVUozoMPpAALQDUjXYIAEHozb+B//5hMpj/UOHChAUZLtRg0EfEhwq5/HNRsaIDjQaVdXwoAA9IkiX/LfrHwOTKlQ6fGLzA8p8pmSUx7fiHk+GefyX+RSHCiQMbDtq07eOyaluKTq1mzLBiRY2aKWqslOATK5CxIaG0KQCrIIEJBwnEffmC6c0bC8pUqMi1DRQ/ZPwgyLPEpxWfYCMM8cqQouZgwrj+rXGmKKERRc7+2fs2JqGtT3+cPfJn2KSUhUP+ZVgo+HMG0gb4zOjEq1MnS/syyMuQJXYW2bSz8FuFsuIXTq8cOBBVSoNwURrmdPi3j1euWAIH7iiokzDJcSvZTMeenbDuAf9udES4kqZ27AkqthjMM1dM/xX/Di3isMEUG22rhlxZtYrfPkt9R1idaqopBvxnCb14GcKo/OhYRZwdHpxihwFH4ANBUCBghhdLVluNDz4oCcykUWSKgCFsEjLsEYNUfOchFXF5xBYjDDLCCFuwMQybbyqgkTEwFnhEs5pAC00h0GQLrBM+/uLnH9hgk62QLI6YUp78ErrIAgESAgAED17pwoFSgANuHllW2eefVv4xJBdjckqoLfIeOuCfiUxy4bqViAApCpO+2GXOhdpjiLs5OZjpH04SmmAlngQlCbmOpljoiT1isuCfROBjYz5OoNkmPwialEcecaoY4b8Ap9JiKqmm+u+pXHLh5Z8WeOGCl/9ZcOVFQ0so+ZWSTihppZVOQMtgCCIVyoKhQmRybKET/znRn4RUVFGhbP95ZB0zFJNRkW6+ufYRbBT5BIx/YhAS0iGa/cwgJJuawQAxqKRSniqP4HeVObb5hwNE/1EBAIMFAMACTsIM0wFZ4olnFS6e8HAvS3gxRjrpIE2onYgoKmk8g8zDrgeSnuO4pEW6M0gOjgcGiQmFYknZpPBMkiBgDlzwlJP6VrkwIdCGYKqVVKtSQ9UApRrBihlKKJYSSniZ+uKpr6ZaWGBfg+0fz0wKB7t+EsLxnRY1ynaaR8Jh5x8wFAHDFh7M/eedbHnAxtrsSHnoXWYTymIb0jpBwxD/ecTYZsoj7uUXglW04YQNBjiYZYKCD074y1deiWeOUKiewSmn1KSa5o1rlsggkFfawKTTswMBUiAIXQgllUx6YCXdUF8IZoW6+McBExZKRKFGCXtBUQZMWYQoTjiZY45/IEjo2XgVomIG/6qa4r9YQ29F6l/HB/ZqS2jNgJ9tjvhHDIM8E+16EhUqkSS9ScLMDmz2/+aeNTIzUd3Itq2KmGEhv+gbSeD1DwMYwhD/sAs/xHAvu4Diec3jAAMY4IeCIQwAApgCG1aRoVywgAVLmMEIgvEP1QTDEr+KxUcM8jqF6IkwGvBBQoaRHY89BAiny9RgviATjnBkJSpRycp2/7eQLf1jEgaZRBP/MUTeZceI8IDHQ1ymEJwAYCF8IAkHOLGIMQqFC1lg0PTa4L54xc8ADASGAeIYBCqgAQ3BaEUwHEgJKrywVwbgxT6Ulb4m0cV9E4RUtFCnohMZpl0CvJZB9EbAiowhEwsJ22Bo85kGdsIQlhBHqfKjjW2wgRmcmAUquTCCQLBgVsvhAwueksJUfXIfKUjBX85HCRbAySBBZIjvBrO67FDkAKLoSOxmWEWWAEEjA1giQ7z4kJEw05oPudlKOLAIDXKACz3IBdCQAUFkLNAg8TOIJBgiGNJAMCFXoB71/jFOgyCjDSSJjUGWZZBC9KIi9UNdi87Grf+ECHQhduPWtAgTApkATB7/WBxsNNSJXLQpFykI5CyYodFcJYISHtILX7THh1xYAqOByQAw/sKLVliiFZSqCe0Gg8yaCFN1/6DpQ2iYMmiApJfJewh3EGCSLTUCJENh5qIMYtNr/uMDBkHJorzJhTu8YQfbmAP1xmk9ryUElwl54zkVwlWDyJMh9JSJOf+Rh5JEYAEa+cFgrNUihWKDkv/wx4sgaZJNXJIh+6wJP+QhuAzwAqPAKGlJgTUsSgDDsClAlpGSJccMKCc1I6CUTqzaEYEZxCE7JQ9TQVadplpzqKUV1OQM8lTswACYK3HDRRRyuztA5w25kB4y2DgdsjL/BALjRCtaGeKZrw0mBqhlkbYAqBFFLkQIJVnWQx/CvoUsDoKIrCdd5ikGwf4jcJFVlmdIM17YnC8XoAVJEB2yEoq4AbXrRe0RUceF0xJkIfAlzO3+AYOFGLEkfpCmfBOSQYOA4CYACIRcmvSsfGokrO9TCD3NqhHhxpdjhhkoihbiipr8QTvuOwJwF3fIebrTINZNiHS967Vk1eY1VONFLKqxg2yaRJn/uLFJchrG7KzFsxYGckJOy4DTHuK1DAGjQV7ykpVwgQus7e8/gCdlkBRhTkOtLUIA8AYBjIALJGDwaLqKzop87Z5lrciZQVLckiDhrXPiQVyFpFCGwCjD/yq633HJ09uO7DbCJFazPZtkz/YVWmi1eVdsSEMFqgViY+iNLwKOx03sOOTIpf0AlB9yPIVc4sr17UiS/3GBNWnnFQsZnoW1/I8t7yAX9aENcZfF5oUsSwxqJgmug6wR0pLHBvH1c0UgEGiF6BoZ7OOXbaAUmF4Z5Gb47QikV1JjhQwVAURmQKN2XNqc7XowA7jdUFnGxZskRAYK2QvHOMLWa17kTQbxohctwIIRFG8VQxsMdSEwYYOQALgc08E1HentPpdkwhU2CLEXxy95UEk28kiBOBIxg3+MoBr/uDhqpzxFjisEwOM2CMgJPieWgTohiHjINAdTgIqonGYj1/+OSo5nAYSslwU5wGwsuMAP0hC3I7ReCcJZolaOeRjmMtmt0NVMvXuOs+klnt4/1tiGEPMr2YERBwtKUAKL31cj9b0Dak0O5G4fnTBugO8Qh7gDGLzcJNkGyRz8+49U1yTsMuE0tf9RdmUEIi4LFA1gDZ4QfqOOM/T7R4kQuBAcYGcFMKduGyQs9XoGPSHI+O0adXvsIxRiFbVagtkZMsTulFz0p5cJfAei8opU8yGy1UgC5l53kEhRITI495x6+RZnBuAfHvgHwGoCARJ4+/Ak0fQ/NoH6mrSh8CzZ976db0/q4+cf4sjO2AXlxdh9nAuNgj3zxS8T0Abq9YQRAUj/fM/FmUEqBxKgnfBX8Y8rDIFoIAn2QoofdYXkfzpvPT6FWLzaQR2AuqZ7sguZKL4FjD4SiL7MQwZkuAI6+AcRwD7Rc71AOZ0BCL/xK4kCOATUQg4AK4leUjJI2TjCsDKF4C8TZIlAGQj+2rsR6DiF4IRQmL9t2Aa/OZKF0LWFuALskC5+eYg3M4gSMcCKSIaHSELE64j6acI2Gww1+0GGYEAGnB4HdMDowzwIyINTY4gcUAiVg7aUIQSDcD0P1A4+SYgzXIjvSBk+YcOSkAG3ExTaIw8XJImb+YI3AJSFyBkr0zQPAL7nCYVtKCeiabHXOIImKbHnEzqoS7FrYrd//3grPZufxEuIKNQIJFiIMVgAyZiuy0uIKlQI4kuIKyS+VdxC4ruCPKDAihBDg7C9awoF+4o3kBC5hwBDDywAAmCI7rgBOKyZMmQIGRy59esIk2mJXXAIGPCJlVAqX6iCISiEQZKSxZG85+s3fFoJdcmOsNEzTFwJKHQGcjQJHnmI5es/E2OJ/TtFLSQ+EpBHEnhFOsiD+QvDkGA1Y9SOFLSvf3BG8vCT8QPGitgihTiBktEOPUQBkEhIQYmEitBDg8A+EiQJFUBGggmqhSAETwOERiiGQBAHMlAfHawLCIAnV9TCK9DCh2gDousI6/HEmiCGtjpHjcDECGguKTSIMf+oSSAsNqeTvIWYMHvMwniyx3qkR1a8As7xgCowCAxgvihgPe2YA5ehIjUcv7tLCPP7h4fUIoUoyNISS5nwyoc4yINMiEsAhIQAhInEgyg4hAzIj1XYN5d8iAUkPEITLpm0piYYDE5kCHVUCCQQxZ/8h+dqvGKjvFOkvFUkPKbUwqZsSTrAx/kjmZR5t+wIhOkASK40iDkUzYU4S5Bwr9IsidMaABzAgloABECIg9nMhkgQAA/aAQswBkIQh/sAmjlgEFAoviAEruhzvuP0v10bkYUAqJ4kiaCUDCQIyoRgR66yp+kbtsd8wHp0SctchaV0SVCggyHwBAJIgPRTgH//2MyEYEbCyJQcGxSTeMg05MqKVM2EqMWHuAP7FEgLawSjYoiyExSZqojXjAPZjE1raIQAQBhMsIAiAAELeIMACIQquIHeHAIEkAs6mAdQEE4SwMs2WCOZAAWGeCt15AznDDIjDLrfsqdhg9Eu3E5WpFEQtVGgsY/PFAD4JKog25L8VEMY2Mj7FEgBuARPq8W0ZIjT5J2JXIlqogCOYc2Q+4daONADjc0FRRgPegODoVBCGADfxEwGwUJ4IjSOcQwV5Z3pjJa3YtGSoIMjkLxtPM4HfEC8bMWl9ELgpANQ2AZCCBQB2IUtkUqWwIP8VEaGkIOIxA7b8wVFTQhGtbCH/+RPIiUJr2xP/6yII8MDJq2JTDWI+hK52JzNA20EGiAEAqiC3kRJfvBQUJg/6gnCVEy4CFsIomsW9oEXMvgHyTDCEy2tTGIIA/oHM7ABXjUIo7sFg6CAKvi1f2CEhKO+36JWGW1A4vtNOpiDPLgCTsABHBAHlyGHLQEAsKwJIF0Il2HLF6DPwfjRfwBSSU1PC6MB9qyZxrym9WuiRzWIM/gJb/M0uEwIHlWmdlUIN/yHRC3LjkCA7yDGf3hLg4gDNIyCWuEHwaoLCdw/s9LLszII4XMSHSwEHCiEbXACgNmGkf0HMojW6fwHlx0Mv3I8VwC+4DsxftIICAAFlxQVvP+8y/zAD/zQQXEQB0/4TEh1jyioJl8YieQziFtcLY3whn+YWo1IyEHlV+wI2I64QEs1iV38B0GwMH8luK2FWJFUCHNNCE9lQyyoiIX9B6BiiTSA2ITwPQB4hkPYBvzYty7kvxKbVXrarSO4gmchAxuggBXIhEwQBmGQggqogAWIgMdjKJi1phpgCFhQCBy4gioBnHb8M8cZgkDYhdINgNLdBTyInR6IAtY1iCgoiPJ0GUk1246AWo2YSCcFiSjtE+wgzdLKWoJD2JrxhkQ1CF/Y2qMlDOUljKqtW92twew4A7L918GYzYcIgACIhF0ghL1VAOCERRzl1vwAUX3EgRv/aIJMgNxmcIYfaAb2NYhmMAgeSQJiVczEfAgzSD/ywFyNoFkPmBKAoS7qgjoxQKumy49nGNTUHVQQaN3WVYGyZFpPcFqGhJ3gXQi4JYzf1Q5PMz+2RL3h1YWIZYg1SAgT7oiAmw5Pw2CNkNt/kNSasAaGwK8wSAgQdtuSYF6GiFIlmOHpgDIKeIZAIIciDoQjDgRCCIdNEAYecQbDXAj5hYVBWIFB+Ie2SYgFeDN34LDB0NyEqAF6EGPM7d8vfohBoAYPSNkjWB8idB9do0K/1NkMUOAGfoEoiOAoiIIzCIRq8gSEBUY3DASR+IfaTS+GMF6vLYkWPjq2HF6SMGEU/34IT/NUk6imerWmZ8AD57WGiPU0PKjdYgCJZ2AIpq2Irk2Ih3Xef6BbAK3aRFaIpyIAtx0JXzA/AUABFKAAd1BH+V2Ic/gHPehfheAwJ+DVsaEGaviHQRjmhLDihfhiM6YHPVDHuPKH9xWGJGhmhkBjHAAVKSnZezk2qpu6yLync648EN2GKiDdQHiBQECBF4hnUL6EMzhDhH3kwXjhwWDkmthaQ+6Imh3bhPhMfySMfH4IFI5kjtnnASQJEFCmM+DdJzUIAFWIVZ6TM0geHtWIif0Hj/6H/0wI6K0Fj9SIgEWBOkhcgwjA+NWDinhmZR6EZx6Ml2YIRYqWZoDcTP+ogcd7vITgMCXYBRQQh1CJwEJYHN2a0+uk1gfEvKdWSYNoEHbm40FGXpM2CBt+CHx9CH9FAWWqXYtW5GvSYPI4SIQu4Y744X/44WswiR02CEwGCbQ2CU/AXVguaYbA57DUCI7esJIQa4WghX+g3o64hNMlbBTAAApIAvl93H9whmagB82l6YRQZmVOiJ9+iGauASgmjAoQZmJ2BSVAAQFQgmfAgCrAAQ8QgfyQwAh86gis1tl+bVKQwCuAVaUQh2dAgQBQghz+B7cF7kJOCEbG7NKC6/hyPYAmDIjm6302uwN9iDigW4EtCebOao1Q4SoyqrUGiZLOayX4B/EWb+3/CGyWeNTkzeUzcIUt0ANg/ocKoIcV8Ol/0GxYqIEamGmSWIEaSAJqBglfTghfFvD4NYhzaAZhoAc0HgQdEEvgJoRCxQEcnINVyIMEyEdGsHDx3fB89PD82AYEIAAMgGezpUq6/gcUr4i8NonhHusXB4mJ7eS6NYg0gIOHcFJYhrmQhBTsronq1ohrYHGSyGuxVGxXUN9/aIYyrgG/WgHI/Qdg1oN16GmG+OkKgO+SiOySkF9frgBnqOItUAhSfgheJUZwrQJfQIGhtuU23wU1R4HP/Mzk2W6NKGyNeNgXJ9s83zV/VVuSqAPykOTp/miPvt6EuPGK/mFY9vGHKG+N/wibLpaJiRRrEl4Isa0DcrAmIH8ISy8JGsjlsDxyzIXcUtcDVxgEYSjw+I7y+M7mFUiCJGB1+E5TNZ0O+K4AKl6B8k7uf5B0hqABfg2Aw07YWgiArI2d8n5zZQx0gxBb3vH0wbBr3sFXPjeIAGBxFu/n0qqDR68ZTjcJo1LGbc8OEJaJ8/7oT38IuZ6T2XTr6fA9GtCBeh31fxAGg0gCJPfsVj9whTgHYM7yKvLyJBiE+W527RDlhBjykqiDg6+IX5eJt4z2+6ymhY8vYiQE8daEIAPpihBphajzkTOq86ZbcGeIhTSIwTYIlI/rOYn2aGf5hZhauUaBLXCFFWhcfP/n94Sw9Yoo8CzveZAAZih+vApYAapMCIcH6r8m7oUohoQ3CE+lgdoNdKXvYBqfkzAARodFrXqNBPAmOA57s+0OOHcwO3RnppDXiJFP94QweYN4rn/Y+H8Y7GyghWxoqo43CFX47n+o119AARrAABwwA4i/6Z0P+IQYesiO4vmdk2ZIAsU9h0xYAR2weJPI64SvhanF6I4g7/GOa+8uCbWH8YqIBFoohlpQfWu4e+PzwHcfDBX2dpao1xOI+eyY/X/Ae7xPiIW8/ZKY2ERniOqGA7pV+YdIhYTg+5KmgV8QzGL9B1lfh3tfCEXikX2vflZ3jDdd9fitgC7necZ3fPj/frwmlvVnjy8diHvUqXvxE292r4i4R4RaYH2jgvrBgASNqOSKyH+A+CdQlcCCBg8iTKhwIcOGDKUIEeJwIsWKEv/RGJjtXzFatQp+RISxokA4E+MsRPkPHTpa2bL9CtfPiRlXApMkWSfs3zqDzv4tIPnvp8CfFYYiRXjuX7OCTZcqXLciSYWjCS86/OWxYLGCtA6KJPlVqMATAscKBARIoDWyCVe4RagkI0lrqtbGVUUwYdh/vwrSjSt48MKwextKQfJPIlaDmUj2JfzPrMFsqjZ+/SgwcsEtbk0qvJaQW6qVv8iIMGPDjMEk/4S5ptgTIRKo/2xLRpgk3Do9Ah///wo8sVtBvBMvCWeIzq3I5v8ALc/dUJBbJMkZht0ovazASwY1S1asuGGDhWskcxMICe1EHZQL9tVEWKXga6oa3b3872vYX+8RPpZbKqpA8g8kceiSRhqp2MCOGX+AsUKAAm1i0E6+HUSUhQdZxVCHggmzwgoduiYFLYFJoVANnhVUWkKW+UXWdRV9VMt7KOG4WUEnpGjQYdsBKVAjQSLEWUEY/MPiQf8Fed52qRRIkg5G/qOYfBW6BY5kbf2jV5S0/EVlQfJJp1IqCuoSDjuK/PPHPzZkUgNCO71WJ0V0CoWhWzUMQpVAOrmyRZQKaeKZkg2J9pUqERzEHkIn/LidaP8MnWAckZeeFVcqqQDiaEOH/uNilwqN51Z5uaXxTxypsCLqP9H8k+qSAjHq4z9h4RmXlv+ABtlBpakiqqil5gZHrwXpIg0ra3TjhCK2/GOLDYrY8A9O3cTGE4cV6VRQT7MlBC64DI27TjjdgCvMOoO4gsGgAklBJplVGuSqQctF965DtZIUlL7PLSfaWukZdAIk7xHM0LwCEYsQQTo0NKFbkwqVcKQUjccDQik2halkq/6TLC4NMeqqxg1TdI29vB6rkKt/PaeqrYS1XBBoa5hkUhrGrlEBGGAcNK0rcBGHUIXrZEtYBeMONlsNuQq0giuuaMLvnHYatBZ9B8H8qyr/TB5kKUVGXrMcShSDTZYwCzNES49pU7QXxQVt7TFCEDP0Q492k5VwyHDoErJDfieU4t4Ciap1rKxIw2tJbq3Mt0DnnQfHGpfzYIMTBkFbUD9TFZQ0hUls4hrTDu2kLuoeXq26QL7txO6IDx3049wFXeyqqHsFXKbMB52iHuK/O8QYRA4V+C+pE0UneUE7YXURrBT9kFB5pzr/jx2NG7SzQMEH/32o4StktYEF8RADjqW5uPX0C70veBy7CoQSKwtpSBH2Bl1f0BoNZMIJ0OqcQP7AJrgsJECs6QU73FQBYXyIITvJyYb+8SGoSTB0dtoJ0qY2iBqkgnwOidxBAseQ/0EpTzCpQIeWckSawaAMeefzGAmH1z075AaHIzOIxoJXPR+e4hTRkJX//kE55xHRiO+7X/A0lpD7/aN6FSFcEhniJJv9o3EEm98/6DeR6v2AUfcjXEMu14A1fGNaCJEWNVZQtIaE4x+9EAgpetELRWDJda05iDAGwRuBYJAwrksCGBxEDXY1gxVQVIgUmiEFHqSCjAe5XzQU+Q+CxcBF/liIq/JXkVXFgT7voqTzUAgJKB7OLcmaCGgW+SsRJgUoUlhAKgsyjYKATyD3syRCjnhFu51HGjib5PBYcQpjloZgrNjhDJtpkJGZ8EysSNWxeoW9XxoENLogXCUbFw07sP9CisL7RwQKdL8qGtGK/xuDagTSOWmZoWhvTOAKzJCMgsxRIA0MAU6ex0drZeKQEgPSOrphhnyQ4h8i+NzQWnSQCHTse6moW/dehQtmmlAgm4Rk9U6pS4I50WqeJMsuGYLOZkgxooKBYjPMF6RV/uMbcLBDFV2py1R48nDY298/HvGOf+AiGsw0yBWxKR2eNoCnRjXIIu1QM4cMVSCNSwMrnjqRW8IqcLpQiVOzWBCbFmSTBUmi98zTgHv8Q4D/CEHUwmEGttIDawmZ5z8yEQInMMIg+cAnO5wQgk1gqTXC8GBsRFdBOyGtG66Y0E5G0Y04CmSO/eiHQFwRV3+AFZc8UuQGFNH5KiwKJKM27eY0S2sQSLhUMEE9SM4ch5AoqZQsQQQS93ApPtd+4x+3LEjjvKmQpqDUQM2AREAAACH5BAUKAP8ALAAAAAD0ARkBQAj/AP8JHEiwoEGDdg4qFLhmYKSFEO/9azgQDsR/cQL8E3Cxo8ePAyVyBEnyX4N/Xzw2TFjSI4EPLWOSlCBT4COD0QyWoHlRnBw/NYMaPENR4EmBLHgKBCC0qUB/Tj2WEkjkHwiB16JG1bhwkkyuKQdeUhhHK8E7UV20RNeSa0cFAkOZLeh2rt27eBVyaUvwaNASebXe8Ihg4KKF9Qwec1gyEqCC4AJXDAxDsuQcWiAm6HhoYCBVtRagUCJwRA8VI1SomBJohwXXO1RYCCTwxRnLF/3iPjh16m6QPCA2G/jNGsEXv3EXJshAIa2BygqmOpizo+7kMh8IBKKwMnaB33YP//jHYsrBcpPKCfTqVH3Hcu7L5Yj1j9K/RALdBE1s8qOu79ip9dEORQgkQQ4dDedUAYYZ9AqABnEz0HVBSdQQhTXZc503SyUHhAUQyZVbfwQBRhIeAy3xDxuhhNJBD178EyNJixF0DCb/VNNRjDzKeNCMBJUDpEGT4AiACn5w8o8pUckAYUkMLNfSWGaNJxOTMbHR1C4QmaPQIxZBFGZTboVnlF1jFvTYQXXtBtdmCmF4UFUHjYTUP+aR1CNIOA60zEJD+igQkIEK9GdB0RkEQCycKFnQSXIKZKKkT37UXKVC1YEpRKgIBJeIBX0BhBoXFVVSIwWVRWJQUm660E0tRf/aEToaCdADCyRNMYMhueSS5z/uGYTJYuVgEqN6hZb0p3YPAMEssP88q0yi//RJkK3jpSIRpAfFEIWrQsn6zwVPNBWBQZ0FdSlE3y4kYEvIFQRqSQj+UxesBekHESsHbbtQZ/gFZiZEdM5FQVBAETSBHBPZA0cqvvwzwj/UHpRnOVPwAYxA2pHUMbCYfExxsNAaFOwUIxjC8UIYF2QefEt5BUAgiPglqwzl/lPGRxwMtC64BzHRF9DgwkUQnBku9IF3HQUAiKlzDRxRRwF/NF1eEuAqQyX/dPDPAFYKdMJESkTxq0fmGTJxtAYpo1053EU7RcvRvVzO2nwUpF4ssfz/qkYwAxnCSy47CDRD4AIFMQQVaJCqELJG7hLZmUS7inRT8yoEdeUFwQOSBIX/U8tA0yiUSMF1cg4RU//oF3ALla4tECWOqyBQnrIT5LhBv+bAx8vQAjH3CMCkMALKKqv8D+BVDCFJE7fcEkwP5u0AuECMK08QFUM0IYkkVAhUBUFVoDFEFv8MccXiwRwvEB+H/8osxoFUUw0Ab+xA2z9XR3Uwbj1bUZz+wS/V2aMmFxiIfVSnlWOwh4FraopSzIKrhdDHdgMxD6lmIDs+5O4fjsDTCFphjDyJ4x+3+McfyOA8SdwiBH0IAUFieIvvSUJ85aMCFQyQvibMMIZ/WBz2/9BgAOelEIUD6cMCYtAEA1RBh/9IwT/URpAZdGIGueiEQiTCkJg4Kjl7GYiStgGSXPyDPvEyiAaCcjkGWoZ1AuFiTYz0jzRNxCoHyQUM4hVAN4LEAQLpwkV0cRuCzEIgYZRYakbAyBEEQ3ljoEAJg5ELS6DBYrEIxC+QEAJ32KAkdvDHJhawxBiYMjj/0EVCdMEKXODCIk0wwzhAAoYQQK8JitiYQDoxsU6E75ftC6Yjn9EEVHYEREGBxkHaUZPmLOJnflzIuTrykH+8AQQlYEICEfZHj0wKLzqC0Ni4hRcneUSQHymBk1pRgAnsZQICOcw/dBCDZ/SgNIawxMYY8f+PGw6hn/+gQhDClyeUGeOIIMEFS36jC3C4Q4iJC+gQ5IG+IRhgoBcNggen8IxfmKoYFnsDRLCkpYOgZSDMjIo8/1EYO35njQKZZVT+c5GqCeRBUemCTKOJnc0NpE08/UcaAmHGf2gsCP/QZUGAodQsIEMg/1ECOSiAgRgs1CPGzCouCjKKgmy1I5GxAxMXZ4AMZOGGO1xIRgXaiWCgLArTaQBbBmKFJ3HrOqcIKkTEZRBcoGogyNQKfQoyFVHEFC/wRJ1BzPmPCSrkpP846f5qksiPANUjsWCCZkGCzqGdhIs5UwiW/lGdXLCADwbg4caUKhClsvYiX9UKTVNJkiv/xOSiuA2Cbt2qBhX0AAWGq2u/DMIkTmzAIIHVa15KV5IzVKcjH2yJnQQCSEyNrSDJ/Uh28RIoEBXILDsNyhcJogpfBMINlBhBWoPwyIEg9bWWcK98AwqSVv4DF/bFb2wDg9SItnYgwMBtgINgAEsEQw3HK0ErWqEzgQg3jv844EXgQAOFHMAsamnVQa4yEMaC5CT4Uq5QRGFYwzZFwzUhZ01mKQuZ5FUhKDrIF+LAnwj/QyLbJUhnC2JY0jjFvCAwRi740AlLHC5v/+ChFJMagq+eIsT/0AM99BBletCjBp8kiAz/YQsbOKEkIhjIDfPCwySn9swGCLAl1KYGlPGB/wV1PVtBEnYQOwD3H+m6y7s+sgcR52W6TelzS5QEzYPk7AIs+AXRPGwQppklpYGxQA+G/I8ZzCC+AvlnUm2QiYLQQyEr+AdULOMKMqP51CkwABoYqYbD2Se6BoHnQdpFkAtr5bgQIYefd1OgGnXEBAZJ4DZbwoGSQoQPCbTPNkUqEGbvhq8DyfOdDBIeOYLEB/+AqWcJUsGOaOoFFgB3IHZBDvjNIBhUyMBTBRKCbigElRUoyDsGYkyh/OApkpFiqvdtAH5bNAWWZDUlipoKaP/muMfFQV6sLRBcx8TZm1pGdMLCOQb/oxIJBAzEQaSfQoPLDQzySLIWogEnxMAo9/9ogMp/0QMn7Wwhi2CSMf4h7kAofJQdmaZATu7Vi2z5Iu6WLUh4qORUDyEFSD960pGeWkuPIBcB6x8i/TCBFlR9IKr6B5fwoha1GFsrtOHwXMRek7jtmiB+sClJNq6vPt6leiBBsVNsbZAGpFxDJ7hDKyjRAj6YkRcdYICsOcEAUwyAEC+IggqM4YQ/aGXeApn3I5yx6yUj/fIZSMHRM5/5FBhiBiygBC9igQJdqLwBUpCD4GcxAcH/owUECMQUpqCCGRijMGu8MN397HAIsa5iJQnbk1ygJLcfxOIYL6pB0qi6ZyIgbJGo5nmCkr839OAJe7jAPrhgxrxNKhZ84IX/+J+QC/HHAhirGDNBKK+QGOgcJKN+/7t5LhD2/2MB6/hH0CWTgf77///+ZwmtwAf7QAlPsAvo8AvugAEEEAsTw0EjgGBq0GYUiEUMMAwmlm1NgXACYXwEcWcHgW0CIYJnJxQ0wXz/4HE44GPrERPH9XX/kGPdNhfAthumwAmLwAGzMAuJYAF4QACjtwuREAAA4AUP4AUxAgABEAkVFgpGcxGFYwEWEAsXgHGVkAv7sAr8kAXysA+WwAeAIzhDNoCtYAgpkAH/0Ab/4ENPAkMhYAN/YAufQAoK8Qn/8AlKtAACYQt3gYZZYFaA+IeFkAEbYwm8UGmtMAOJSIaKOAMO/xgMncBvKZALkyUQGiAKa0SC/8Ag1rAGcOALENcSHJZd3wQ0Hgc71tQhlVOEBYEHZCdGfbQInEBn31GDH3E/MuECTLIIiyAHLwAAAFANh0AJHgSBjsMCsVAFubAN0LAKTqgACRCNCTAHuXA/95M/qkGFVliFT1ACRLANzLAKvMCIsXBp/7ANaGgQeRBqTvEO2HATkOdV2DAQ8/gI3cAOivAJn/AH8/gP2PAO/jCP92gLMRAe/dgSvdARWXAE/1AI/0BR25AFhZAFEbkNwJBP+zBR8nAEC7mQR8CREfmH2yAOhYMcDqBTpSAKpTAOJFYKCpAIGHcBEvAaU2AM4mAJvv8SOgOxZwOhkzxViWzAkzJhLRcBWXOhEXgQY9qlEEi2QAJROD75G3AUExwwHpjwBvgDjFNwhmiYjlGUWlTQVsEQCIzEQZa2YJSQlqJniIYofm3JC2pJCfmUAfzQkOn4hwJBRrsBFaNmEDcBZQKxXwMheaL2D/FoF/JAEAxJEGooBkewhQagMpSQAvKwCsiADB8pjjswBTuwAwDQA9CQDq8wmulAB+mwCpwgDpTQCkOWlp3QCrygDQWIk4HwXcamJeMVFDjVEWwwWkIRlb/xASE3g7/BBdtQVBwWlYw1bCDhcRchbQYBaARRADlTiQqhk7vAFGTJAloQC/twBJqWaQf/kQFD4JXrFhNq6JAlmBdZBhIMKQYFoYZtAAHr1gZPVZcCAQEQoIaXKQb4mZj/gD5klJiF0IVl9ZhHsA28YIjKNyBWAZxR4Zx5YZ2viGTgkgZB4ZO4Mlj/wGh6cReXZRdLgCu2IwBY4AGhkAcOeT4LgT4fmYYDAQEXwZ/rBqDryTkyehAkABLyeQRP9ZFAegRtIAbIMASFQDhT+RGviB25eaMF8T8K4RYutRC0phD3RFkHMQdBUStRAYIe4QEeQBCccAPjYxfwaRmbEBV6KBlIACA7OhAkoJ/IsJ/02Qb2iQwkUAUCEABbJxBcQnEFISXOFopOClwoUEgiRiVRYZ0e/4EcjtYS0hd9BFGlQXGlH6FwBhEHj+EWImUBxlAF27AKdAAKoEACphqnqAoBcbqfbeCjHymRC7GYBtGmB7GmJMF+rtCe+ycQOmd/tuoUdnqeIPGmBEGspfoPJFCqypqszGqqeZAH8QAX34KCA9Gnv8ERvmCtfmSUEVMpafIc/+ClBeELAdCtBXFPd9ADUXAGiCoUYQoSIPUPjWAceACoBqEDA8EwEKGtMxeDMjFXAgAAAoAHAIAHe3oJWPABBEAAN0AE4kAEBOAJ5PAM6gMKELAK/4CZV3AEtnUF2+AEOOAENmADK7ACW1ADmrAJFbCm+Qc0sCAQ7DgQ6LMQV0AC+f+wo/M5p8iwCvp5sT2bqkB7qnlAAkM7tKWaB6BAB0q7CjhACDjwriWhESH6pAJBAygyFnigrXNBAB2BBcihlARhruGKR0GlKlnHXDFRDEMoEPG6dUv6D2NRYbjxEI9BC3/FJgdBCFD6UxfxtjJRTeA6EHsrEL7gC7Vgrp7gCWHQBOGgCf9QAfH2D+wHuTUQswWRDP1ADaUWFFZ2DgOhIM2gIHpAZf9guQLxsv0QCoXwkY6JDGeasf/wuoyZsaUqCeO2C7uQtbtwBlfBYe1KEDAhuAJxCX3Ktf8AtcdLEH6rEBjgpH6qqCBxXbWhV4AACFlhEBgqEKpytwWBryARBv//oGsgMbgGwb0dIbckIa4tkXWoYg3m6xGKpqjeKxBYcAM3YAZb8LgV0Ax6UAF6UAOukAQFEW+QWwFJULk1UAProAfNELkL4bkGYX8EAcGPC2pbwCUgGAZhgAE4cAV5kADPmgerEKc827Oqqqo1e8JxKsJXIA7iC730CxGKdhCYOhDzaxAgVQzGYRCKGxNmcBc1fBGjExhDLBBBDBHuABHS2xLRkL3ZW0cFYUeBaxCqcBGkIQgk0bz/sMQCkQ0EwRZVXBJCUBDxqhVPXBJcTBBFLBBKgAPJ4ARO4Ao1IAwDTBAOnKYCQccHEW9S8A+eG28SLBQVsAJzXAEUsAWIQBAs/wizIDE6Q4yv6lsLifwPpKEEWMzG4DrFAzEIF7HEjfAc4BpB99oSm/sPtOoRl+wRP5fGLaHJAyEaHREOwksQUiC9tnrKmKIKYfwPkDAQBaQQtWwQkywTgMAW6CDKBrEGBjcQdcurBuG4WiEN2msQBZQG9/hlimAG4dBp+jcX+afHF+HABIHLByEMg2y5dOwKfTwQ5LwQc6UQ76doibzLAzHGeqiH9NwS81wT7/wRN0xeMVEDB8HKAqEK19sS+fwPipbQMqEg/+DQrjJbcPBKrFBvA3FvBYHRA0HAAqHR0iEQ3MDQNTFb/yDSdfwP8icQafBVPhXFE8EDTgAGBPEHjv/3D2Yg0PuXBPvnbt3QDWZguiCRBOCsFcKwDkP9D0UtEJz8D64gDBGQ0jFRxdMRHMGRCiQNEarADVJnNaqw1QZxCh6dKloB1QZx1E2xzgoNVf9wVZLxl+ByHeER133VSnn1y1DMLy92bz/wYvN4Cq601hj6H3Gw1Wi7EEfBXNFAU9IcB7oQDY/wXDIBB2NyIZTzDQ2wDopQ0+xmA64QagIcE3+QDASRD71ghwPBCOGwCS2L1KwtDADsCp22Dp/tEUkg28Iw2wKRBCvADqL9D8nQC3DcDwm8Aur8D8GRVxZt3AOx1boAB/zyH7ggDbHFCqzQywTkDwXECnZg1xeB0a7/JN0DQVNnLFQ5YRHS/BE/ENYewd2+zAPBgdEQXZj/IA0F9FxpIN4CYUz8wgO/DNkE0dgD8VVsfdHNoN5BMeClIhCN8BDSdxFMkXV/yyEcMrXnup5lYXYFcd4t8Skt0dJz0UYDEUJC0RCFLRDRcBsmoiIgIXxPwoIqJhCMZhGf5bwdUV0fsQgsHhgPccbIjBdTeqPLLBNv8g8gPiKUU2cLIUcsoaXYscyOFRU2LhOVJRBeUxJlEeQd8S47ZhAMdxea+A8OMBiEwVLMsRDK4GvhUhANHhNJ+uRaIeJBBZ1O0QFeU1SpUQ7hNHIg0SPpURDhdDvkQRCw1hT8cR0vJxAU/3fV/yBrEso5POHhFyFh/wAE3/UkvhkVX3TpHxFBByQugKAbogyMdwTpJSHN3NLPF2Em2iHiofURYGsXihpyUREKh2A7x/IRer4jA5HrC7EMwaIMLGBGaicQndIS3lEGhx5NctcRy9sSQECthj0Qkl4SCZQIjV4pkXANynxjWiFHWK4SqA4RDZFjMcEdQKACFF7kQ1MQOWAieTbsbOsNRTwCfNACEkAyLVEjQrLrf34RMeIVvE4Qh1IQvj4juAgAIHAITRoU5I4p1w4hl4K8N1rsCpESGD4Qu+xT0E4QcXC3ARAAcRAe3/4RaeDKAGIR0/5hNZENdlI4gx4khnI7fv8XH4jiBe4BJMew74eiDAMPETZvPwCwdQLAER//8RzBJUOf9EO/EUy/CwTgAYUhmAdB1n4mLhfABMSJKVywLguPF4pVEE8YE15MOT+OgieBoW1C6jIx8h5RFbKOHV7dNG/AAlcqMryjHVMAOMDAqANh93NRDh0DH/huMgehI3AEAFFQBdb94gMBCbSW7BZQ6XehxdHE+N/BNRehbTUR9h+RA/WCGxgi5zIhnQQh1+vpNR2ABdwwDXDwC1FQQX5vMbvyD3z/Ee6BCeWQKA9QexiEJ9BBENoxc5c0AiTTMcFASTMgZwoRTrUwMOISWkxgO/Z6EJqOGyvVEYKWM80OEdH/IAjBWxDXT+NBofYXAVRFwfYHIS4WsTkQrhC0uBC9DxFb/hG4kgiUUAnposVYsMX8AxDkVFj4V9DgQWX/gPxLOCLXiH/lDD44ODFij3/BplQMZolXsIpTpqAxFCzQm0BoKlJJkSLYSypogo0wZOifyiFDqFQxNoJiwZ8RhXqp9u/XmoINKi4t+ITp04KLoE6lOpVD1YKesBbUsLUqqqpIvVYs8I/SWLRLX6X9VwuOWLZx5bK1A9VpQT9ss801uOBfiRIFW/zjBfGfmn8qDCJWoRjx0oVa/jn6N4VPjoqG/zWR9K+K538GhhQaoqjgn39/hvTkY7MgFYOwqUhSNOSf/yIwYGz/g10QDZUhZG4Z7MNZEkianQxYGiGxYMIHUzQfHFOX70EG19Oyubr1AlUNB7SPJ18erVKl08wfBFGeSNiCcSJFeupm/foWXAqqGfH43zNjEpsiGNc2UmMKxKaY4bPhtoLin2QgZISRIYaz0KAQ/smwDw07JEMSJ65g5IorPpmKkRAWaAIYYI5IoaAg/oFoo1b+CcIAz1KgYoRddPlHqR+pksAgHyu6io1/kKyqq+tMKSi7+9KaI8qlFBtvAqq6oDItLwD4B45/4IILKi1geCqPgsZky5uC6COvnn9+qMiBfxzQki8u8iTnFnHEAYaXPzMopCDbDAGmoFyQQ/+wsh7IAecfO3goEi3rDsJFF1b+wcWgTFmxo1KsYlggBh4WIONQG3uzsSXeYgTGAJdGQMFHIOVSEqoX/glFFB/uc3JLrKCZi5B/EpnKzYOYYAqsgsQD9llooyXPBLZk+Oe7g/RjAEtdzjCID0turIgEQg+6goyCRpjCmCo47AarTaN9lwdw3JEE1YJSyALHpYLwNwgqglB3BCXEakAVggqywiA8qHLh16dWQQuuWg/iRFq2xmGSKfS8sqOR9cysahwHxsH4ZKwwSOsLlOfy9pd/+IjZkkNrlite7Tb10cdKJz0IVB5wYaXUg1Tt10YcDbiRCgMCnkHdHlD4RpVcK6L/7J9s1Gx5a2APKfZrg9TbWpR/TDa5vKug9KqEN9IME0yD7ItLzqXUZusYtMpQ1qCK66yq1kcuWWqAfy6G+B8sdPElilximcEAHF+1JLR/Do0xxoLw5RraGztv2pKZpIvliRmmumcpDthw8uKDrNx8c2dfn2qZqcgmezwE4vruiaqpkhtlLwoSXPaC9q6EKdb/OaGgQGJuxRIDWplBJYNSiDwFcSQh4B8K/gnnn+zBr/wp0wrK1HymQNW05VdvfFVyYGZSQ4UlzpKRLSkMsiCKpWK/zoUN/EM/Y5HZ1uBEnoXNBVmqiNbqqnKHuzwFEMTjS9/+0TumtKMgpTAPLWhw/4ldBCIXM2CBQSZXrspJYgv+gJM/nkKPiqAGQzNkShOWogc9/AOGBdnhP2pwA96sB3JDJCLkDNGfETgEWwVhIFoStjlyRHAPTfmHCygIFWtQ6RjHoB3LqnK7dE3lBe2Ry+n+EYt/POE7F7BWy853n3vEwUvrKaFXyPgPCwQiEFWIRRINwYvqVe4GmihIEnrIlEeUB2cFcYVBVmAGcYznRfkqCKyGaD3IDQFyM7FCEs+CEWuoiVgFwcD2toAxK2JlidpJ3hUrogAwPqUI/2CZF9kyRSrx4TvHM8gsXTmxf5zudBasSq+Yco8GJDMGLxBZ8aZShwuqIAp5pMEYcFCQGP/wJZHvOIUwoBUB7ezmHy+ynibLaUnrWW9HM8hBLijBgl1UhAIDHMxgKgIzYKXyH4iIVgDnAoK2/fJZrdxKjf7ByzYG9ILRKsIOfCmXNHwjSsmk6Al6oMt9nKWOBmGAVEwxAGO8YJoYKQgSppLNf4BzKu9gil8EShVyDqElKZBpS2raEkM8jRK8QONBFiAHLkwgqBMgaprWQAMC9OCJVLrVyZoKLQFUpHQVwQR5cleeRehzK2U5SyVkYCWFrmcW4zncejb2j0c04BtrsMMadDA6SuwjZiXgQwlasA9maIsDAyCESC1AiG0wohsuLQhh2YINqoBTsVBBaVoysQm22Eb/nBlIAWUtW1nMUjYFQQhG6RIRCxCkogFraIAQ/JDXWXAhFwcSCYIQNAOniEIDGtQgeZoIFWlwzZgvLUKulsoUqWylmeSJYFmY8oLedeeKpuAOA4L6gS8EIAD/AMQE/+Gl4FFlLVPZgQUUdAFKXCAXzFhFBibHhxmk16AF4QUlStAK+BoCTWMxLHmM8AlSQCW/JioIfvlrkP9eJwMZyMIQBpwFAg+YwAYwRCt4YQiZoVdm0ktvCdI7ghl0Ug0zCAYfYmEM/XDwH8Y05nYrYo9/3HY8xjpIbX1wgLNuBSyiqG2UFNqw9bhuKjjAILQKSCVqrYd/BXHSIprbARUIIBD2/0tiKzrBgnJ4YRLHCEAjUICDUChAAQngcpD/QYA3YMICbcNEY9KYiwtcoBWkywU/VrGNQmSAHxmQXiv40FlLDGEb/zjCPwZFpW3+g6VMQaw/sLEJRfA3BNjY1DdcyI7ypWZ9bMkCVipdkCxkWlADfjAlUtAKNMC3FQ12cmUPPGCaZoALO2heQW4nYg0MIw8dqEQBLqACEHRXfy892Q54XZHp0tLX2snFQZcy7K1Q4i50GguLC1KNHSC7KhBjwF5jgQkAZNsCDwaGjp6WxA3zxwoz4A8LcsELLuyDE41LogoCMYVAqIAP7hRvASiRCD9wgRfubEUu4MsHHGXgIAL/x/+eC5KPrSXyH4hlKWIr8ggXGmRTizzICrQzqD9fms9H4DjHdWQIufLjCCJHhhjEwPFtbIMfn8l2D1xgJ1E4IObjEIUoZBGKXORiDy0A5Lz5wAtLxCLeBnnqU4F1MaPHRdoniyoFfztsGdj6WjFr2R2jWlW+vMFL2QaACkawjzlj5UWUlemA95GBs+9jCPvIwjYysA15IKMN/4DAP5Bh94NkWuO/TovDtySGp9y9IHLnxz/MmwtLUMISnUi8JdzZiVwYwt/o7XCHDUEFgfdZHgi2ROf37U5ebNQgnLiKcltGUJS18SBN57tBPlCQtoW1Iqvcit2WYjuLzQVbivntUmT//w+MsCAHOQACAHbAhW3khODlqXtF+uzKszEl4lBhx0EaO5UxrGfucx8LuQrSBu4X5Pl8lkfHR34EZBwhA+hmwdL/cdWK+PoN7i9PduDfer5j6R/xNMgbfo8WwoGK+UKZa/oHr1mKISuIIWEKD7gCEUCGQdm7qSAB78O/f+AQgTql15k7uZO7I2gDMQDB9LuCYpujgrgjqOA/C5SLVltBufi/tCjA60CW15FBqPCFJhgCiUm/img+Fzwpr6iv8Qg/7ahAI6RAJCQBCFBCCECGVQAFLlABjFBBtqDCggiQf7CPUJCY18Exr0CBggBDXgOTaDAIuKGKphsehpkKK9yK/zt4lniigfHwlrGIgzgAhGDLtjcoAgvAAwEAAQIgADkQh0EcxBsgBEKgABzQM21YBQgABQpcQkmEgDbgwYoohLrTwK0xg4LgxKfIvuyrCsiqCO7zwX+oQIPwQXJJQhLIAyR0RUiExVYEhTzIg3yIh3gwCBFIi+0ZizaMFnX4wS3JIjU8wYMItqfIFf4JBBTki35Yil7snlGqCGsAmYP4xapQw6iqGpJiizjAmqWYrum6BHIAHwQQgQR4hVpcBRK4goJowiZchT7TgwpwBoNohn/AR3z8hwrgR3pYAVioiFAknkaqCMAzyH8oxX8AhX+4hQDYBYiMp0Awhg8gACLggv8hwEgEGAIE6BOPxMhriqRI+ocz2AUB2AVknMGKeL2lEJxifBYZDAVhxIKCoEmDsAHzSAOqyK1rWIpawEaq+Iyp6EUg8opikBYdmItvbBO2qIWlUAIw1IEzIAQcwAEK6MdmqAAYsrh/GASDoIZ/oAaurIoVqIEaEAY92EevoJuKOAd6qAGv9Mp/cAVBQIFn0MErSL+SA8FKpER4fEe6ozslpLt0WAVxCKFAOAMQOAMlOAMUQIFL8AXQQJyWTAsyosOnoEG2KEqqEBynrAqtYAobNI/l2Rq/iIM0WEqqGC1h9AoGogWoUM2lKEeDKAbJHIvu+QdN5AshKIikxAoKoAD/M1iBFXCFfhjOguhHplDOgzgHg7DHtFDLrTiHJPChLaAAHfjMfwiDggiD3FwKCogkGggAp3TKozzPYgDD5vGWMZDDf7jNpYAmGoDNgqCFl0SLbGiE/PyHRuhNJbjB95QL7YQKcuBO7agFyexN8oDPp+BMYIGLaAATOJhQMNGailAxgyjNf4iBVIAKBa0IGjAptLgGVQCEbDBRrIADnzGs5dkLBsqGX8Cn8tBJnfSKNOjQf6AFWkCHEGCH6nOCFXiXqWDOp/AmIzWIfuxHbxqPdTAIb+LKCsiEFUACfqoIQdjNg1CZf0AHFXNK+jyIE1geGX2KpKxSJuILdKCuihDC/xRrzQydii8tCBy9LQ3VUKpIhQiAhB+AhKXIH+Yk0gpCC5+R06qQTqOoiA+tCj41iJ4c1IfDilRIU6aIAFWIgVOIi0w5w4IoQ605Q13QhXBghz+Qodswg3DohhrwoX+oTrRo0qoA1OTkRyRd0n+g1YpQTmGoAVdYUnpYhyRIAlcQy/wpUqhIUww9UyYy02N9ChzdijxNsUWlimGN1oKwLuuLC0k1iGEd1t/MhK3gBqqwU4P4xmyND4OI1jidCzlxIXaluK1ZA1aQBjuAA4WbtJT6Bz79AR6wlH9ghR/QR6r4gQ4F16XQ1KVQCmTa1H7NLR8BVx9RzdzyCh6I2ILQhf8JrQggGa01EJt/+IZwcIKl+AMnGARvXdV/EFKmqIHqy6+DY4Q/GEWsEAZh6AYz6AZbfQpX/YecJVaDqAEnSIZe6AUzcIVMcIUV+IE3MtSDyBRwVc1JGVRHjYB9PYg5nYpmGNZ/uNRU6FBWYIWHPQhdUM2hSYXzkQZw5YYaHVeVcoYKwFrzkAJn8IthbdY3mpRH0YWpvdSDACdu4Fo42JQ36tetqEcRJQ/1mQpiiguKgQMUAIIXmCW8GVeDYL3hyaKqWMDWTNx/+IBpDJOxYBYFGAtIgBMLZYqURIvQrAjaCdSkOIgyrAjV89B/6AAK+s/WvQe4CYx/wIyfkKit0dz/62C2pbiTl9LMpZiEg+BYrGCTgmDefzBe5R0P0TsI4IUKDwgur5DN2J2L0HXT8oje3/yHMpALLY0W+JMDqCgh3T3YsXjdrYgxjKkxC4yE092LpSjdqTjdAPDCNAASe+jJ8sBc7dCqrVjWqWiE010P3/UK1rPA9U0MXgvAg9CBxLWWZlqIb6wVFPPegxDe62CAAcDe+5iuSLDWDX4W4+Xg9TBBqpBJpjAWrznAZAqS/dtdFciBxhAAO/QFAQCAHhaAAEiDNMBfFS7itHBfI34KEaYK2jkG5DWItMWKEr4PL3zDirDGJEaL9zAutOherKDdRHADY3C3ovCSSWBhoTCI/+waixNKQKQ8GRFz0zWwVggmng3wYGlJCCkz1+j1igaYoAT2im5EGTcYLl7rRfNQgdUFljVmConwgoToqSVIozdp3YoY34LwQkd9P4MYIPzzwri4BpZZCAnosZbxJ/Ioq7io3qkQgAYuiBPGiinwGi5+CvWgY6gwo0iwJcnYigUG5a1wYay4BB3jpfGAhrxIY74oiqpwjrSgnXKQt3/IuQjSjsAIjPGd5NbzZLSgBSAh4ql4KMzAClb2Cg44EqboCvkdiyWei3JuGWD2CjP6B1+6mrSIZ+1QigXmi1WChkOwgEauimp4YuIJnkkoM6eABtRLi+21QG62o/u4v6rYZ/+2GKskOQgteZB/WGdpkU1OwWevQApwTouO2ZxxlgvN1eb3gGGo2N+GGb6C4AJCSAguKQrnCIBsK4dJYGascOaDcGaargifhoqu4wIkYR0CrgoYKIHxbehfsz2uURtVhgqopiBm8YC0mCCtAemDmOeneGftAOIU9orw3YpXZgovpt6xeI+KeJQ8LIjA8I/rkIiEwLqDCOilwOugHouh/oczBgA3eGiOoQplET1czmLzkIp2FsZQAAtmuV+DHWxLdtNy/bW+sQOuxopBxoqEiLJyoB28/odG3jqDAIAn5umCiLKlSIiBpuk1Dh68geTsKge8OeiCmCNXLjZO5put0N3/B3YltdE/FV5otCDutAgFfXrsipgGj4aKkUZDjL2PNUiDwx4PN54og4jlf5he9v2HYNuFHthspmjk/sgFmVnkux7vof7s1G5m0VaGcqDtosC6H/ZhV0bJAIiEYmgEa/WRNEAB9M3aye6bX7ju1lwDr34Kp2jGtHgB8XbT9gDp0FVug6hug7Dcg1gDOuzGhYju5vbc9QBrrknrKFGFABAAC4iFjdiKcoAIYMiFFrSI0L6PvVbmn36AcngAZVgGiUBtWjoERH5nTEZsC1xs4hFmtkBYksxCpqBYuBBHg3huIscYE++BElpxrDCMAJGIoFjtp5jxsZiCFleXvq6In9iI/6BA7R0ghzEVqPKd8pNBZb6g8H8g8aXIAckogjcIgKNcD4qhkrOmiqCmvV+i3X+YAEP/B51cA3QIBBX3inJ4cLSohqgCgPg2iM62caFIiI249JqYjoPAsKfA8qUAAVpAio4p5zb6AqDkKL5bot9GGX3eEo4WqA+4gzvIbGnxBl0vCImScq75BR2DitFdAxTogWE38/jjg06IBfej66fo8hynaYqYNzG/dKEA9YwoiMszDOcoBzUACUNgsOYoc6bwhboo6aeIdVraBQwnnlsx7qeYXretCjtI3akgpO6+DzqPiynhi6wBa2Dfkt6L7mP8Yqog9fEQi8CQgSfQbRrQAf8zRStpUAJQ73CoQAw0oghlUPiICOpyGJDpcOYTMggxlw4Ia7UBIQnfWI4R2IEAAYmYsQnYSAGSgIguNwiJuPRqeIO9eOe9gfN9N4jdQguZFGYkb007x4oiiKeAn4tArogDciU36IBEjxIvgwoNFa8RUAEWYIGHt4RDEIdAQIFAkPSD2IiFoIgcaAWRcOQW7/R/KJ2ZOAhDyR6eAIrKkPmZ2IVnYPmCqAIqKLBDoXk0oB40qIJXuQVJaJqZoAyKiA69Lwf47vldQAdd+BQ44IFU2OS5UBsGJ49zLgjjboDArWWhp5J6n4oOP0qwTvCtEPEtQRZD/ocARxkB3odOKIj/k36KBOllk1cIhkgMPpDrf4gOLKyCEZB516AC4Li73WgCY3i35T8IoSyaIbChHIQN6gkiNJCE3fiDW+AMYDiif3D0YnONyM/xwygIVmOefxiDtzAIzGUCp56KaRxQYKnqHwEIVv+e/PuXqyDChAoXMmzokOG9hxIvLDSFENo/DRI3cuQIpyPIkCJHJsxG0mGRkw1R/CvxrwxCLrxyqWmoZsQ/NVNy8kToCGG5fyz+7Sxn7F+TfyH+SKryT9KQJk369Cl4y5YtMMiGIAzyj8pXNFWqGEgh6datf1QlSfqHpiAVNFAVNQmRtmCfEFANGUJDpWwwnAlHTDFmqNXCjyod/8oJKeokA07/JG8soNDlYolzCibI7Plz5gYq0f2rJnFNHBCgVw9N2Hg1SZgMc41Qo0JNjoJTePESvHOGYCAIlU2J9a9K0rv/CnH994dhn1tLFUEdMgQqW6nQ0xoAVoUKsEJk2v5T3m0MOF12eJD9nqL5vxk8R/hNGEzcvzQJRTPELJHDP2wgBCAiDGmgEUPCiMTAPwDC5lkXD4a0gQuwOeDZGqLxJxJpQT2kGGgEjGRNJAiV2NAhEp40QUxccJFLLDWpUZMNYzxT2xTBdEIFTjshNEVhY6j11EhO2EIVVWr10c2SfYyyyQL/8BADlf9ckRAoCrFT0Arh/ANFQVxdh//QW0TxYck/BpRV0AiBjfGLQN8s5uA/i1i02IYgAcigiidd2Oc/FgC6UISDgqQMQh/l6VkNnp1YIgCGFqoSF7O4yMsQwAADniWWUGHdP2PcEJghaBoyQiA+6jSCMej9YwdChfyzTUi4SFmQLv/ogosdAiFka0ibhLqAO3aRsek/QaARjCFgAZNCQWh+9ZUBz+jSwBpz1pkQZQqF8tg/7azGp6HlbhQHQxQVVIm57apY02cauuvQpCGpO4tCA+iwwI0+BnNQQUmRBxcfBc2okzEs/RNlQTEoBCtDuS4mxELPISQxD7rwsEBbYIEVRBB/ZZCmAf9kkEIQhgA5AsUFZXv/0iIJcdAtQq1JaBG58ypEZ0GlPFiiAAoxoTPRCwXN0BsOqbCavIP655kn/wyNEAM488kiOM8Yh5MhQQBTEDKM/KPIECV/XQh+CN3kVFUMQbwQsOWOwYMdCzQBbUIGZDDytF6B/BcVM0yBqsT/fFOMoD51JCDN3iYk7kMvb3QnAzl/BrlKj9ULGwtllDG1ij4X9GfRHak2KCT/RFRQRICcyJEEpYPOYuX/MMhFQWkEctAIM6BpAFgFfb3cP8jgXdAY5PxjTCDHjbGAMwvw4FCuhZeriy6//DP8PylkUXKyaXYF8t9BBFbYL/yhk/hPpSO0aEEIFA2/SvQ/lEYjgKbI/1ApF4o+r/1KRwiRHO0Y7iPJLggBHD6oSSHBS4imvlII5eBKRbay3kPixgr1gKMJZBjCyeCSEK8UBGQlM+Hf0LAqcuiHNAqZAqIOWLQDfGYcG0ldQiyTIh1Mo2iy+IfPbCghnr3GIUv4hxVKhwBCnEKGgCJXLdyAGD4A44QK4Z4IORK3z1SPbg+ZXkFYsR4iJQt4HTFAENBIPjQQJhBRoEExGPKAggCiITFzIh4ZAi6H4PAfRPhHivbXQ5DgTkL/g00hNwK6f+zCISyAgUq2CBpMxBAki2SIEP9BuoTY4x+iWZ1DYsYAFmFBYrmYAQNLhiYsOuSB7XrbRtKTGTTSMv+NKQPSFHoQBRYAB4kQcYiAEnKGpf2jM3l0F+Y2coKQ4OEzmOjIIYsmm3+AQD+S88z/tvCglJAEBjp4SDQRAkp76MANC8kZnVJxiUC44ZSWOCEVANcXYKCJhNvrSkIGJhJc+Go1+lRJLWl5qinYJhcXcMnTRgJLQFXojg4hCMAUgoqOBPCYFl1NwV7SEYL8w5ylC0DiJJTJkeyhIAAS0J0QYoEenLJUJQsGGrqDEPAh5GsR3KeufNVPi/otoFXs1AgIM4JWlLQhoFRIzO7YgGhQ0yE09AyFRlIJPqhgfxypqEjqcdGHaGCPniGX5UTCHxCdpAteDYk03AWPf5yVI8b/CYkFBNWKWFiCF/JpRclKBq3uKAEXp4jGIwL7CFzg4gfOyMQKbGADMogDPghRhEQkOS8rnlBNtFRTGjthDIKqoRUHlc9JyNqnDfzDBSlFyDcWVdStsjYhohhHW08CIIduJAqZOR2hStGFCylIJUfbyBfqWJAGiGYNkfiCRBCkkLNiVSGCYAgImpcLPhgiPv+QFkIyFQ5nPCIh79CDQuiBkBqYASEhMG9CbLERMyShBu6FxQpc4YqEpG0hrDxjQSyr3zSiMahqsAIfKIGZHYyErJuDjQs4Ib/WthZdRKNtRy6pun88ohGXwCMLkuiQFzjkmgm5FkOSSZJgbtgCBh3K/wx89w/4pMAAksBAMx7RjAokBLwLEa9EzssRGzOkBvNVkX6DrCYqBONgrWCXSmhgAdse0LYUKepqWcsiPzREAMjNzDEMCAADIkREDuFE8xqiroLgNiFVK8hpHXIHhCDGfakA1D3quAzhcOTAsHmBBQJBCICNoBO8uKIkNNGRHywmKQlpVENqgINBCbksaqIncG4S4H/04B/WWIOH3Ufa0v5j0Q+xzFaba6gsd0QU8nvmoPSDkDEvJGnmwsBORQLJjfz2H3QmWiBUgOcooEBrwDEEprpXsiEUwgz9eMg7zDU9QT/oeNBqMbQdHe0UnOomI6DEHip9DUxf1AUkNhQGRv/iA4bUAoMjOaJDFLCRLHP5H0xt7UGQ/ExXzysiR1UIRznS3YJ0kiMaGbdD7kHcBvCAwyLpgQXwHIhdjCEWxsgFMpxgMY44rCDYWAihATW9ivMAjJ+ZtrSlzYtWBNUKnaAEC5CLLdiIoF1I/sxEVUJvGaZEGcuIVEMqtJEow4YJL2/JQgw+AIRQmcEPMY1InPC+1BL3F1FIaCJYhBASR+0FulZBIJ6h9I1EQCLJPub0zN2RaacA5C0GRopzkAtKMPLNcgLkP6jshwnQvQOEcDAtFPYgyQhI54CqhUK+LRERI6TMJyEwaJZxZZX8HJgOYpwiFSKDfyB+IQCSutH71AD/pjcgAj2IhX9KAOqEODS6LwiEVbuuENUjhPUb2XdBIFHxL1q07La/ve3LZgA+AIcSiXjrhE9AhFnQvQV0n0AH/pHWfyDC8BKqUOMMVSG/O4TwZPZM5TMPmogWbfLczAwiciXqhihXIQ0QOHFPwAI+sIsS+wD+PyyyCA6wYQJ3WLIKjEGrgkiBIYYFydchBOxpn0I8G+4dYNkZQu9ZQiyggPg1gBTIwShxwfFNgB8kDCEEQu80D4JYH9GM3sFRWkEQU9Fw09NMAaoRYEEUXUM8AbsAzOS9QeUxGSLZjoPYTPb9R0EwwNCFxCSIRLZs3vk1gA7AQIDtQ8Fc2z9YCr7Y/44pDIAxnJ4KRMGiMcxDOINEZEJBdNcALsxCuJ5CzN4BnQwZvkcKlOHJpACRzQAlUMITgMC1ZMgCiMM+uMgEWEoiqAAuOcIUzADwQc5TrcYHqOBqAIFgEGJBmNamMQALLsQhFgTbqeAELMIiMACAJFKf0MA/pAIt7EIAKMETXMAF7AMlGEfBuEQu8AIncAAHDMD9BUIsvIgTeJoVLgQWwgYYMoTH6czI9OIZgtAvomEQtAIftEApogArNAAcwIEQDMA+JIJ81IZOTCNBzUAu4M4eAdxiCB4ifkYRPOJIfN9DSN0oKUQKbphEcKNC5EZtGdwh5JtDmEC7JJUpVA7def9UAORPI7hOpFTDD6oECOxAQLLABexBK7SANuyDIQTDPxRMGaTYDCBGLPABKRJjMGTAlSBE/93iP+RiLXqGetkAGHwCQ5ACSfYCKaQkKRQESQ7K3uzNEGQBCL1kBlhCK7QCb/ACJcDIW81ACaRYUC1BbUhjNT4BAsgCuATiafDbZ7xcJCaENoIERqCCujkVbNTaZwBB7FhAMyFVQvTgRoSUZ4CjQrjaCxhc/G2L+9jWANwJG3DAKDHAIXxBAARAJADCPp7IHCVE/hSEuk1KWyGeBUwBH1yAG+ZCIqzCKvBDBlABHxhHm/EBL3QCH/ABMXaCARxBHoBEBHwkaBjBP6z/ZEK05D/kwz98Akl+AimgpITwDUK8ZBZkQGzOphqeSScURCugUkTq5k/+JHCkWBBYgjgYQhQsGFuVX0M0wJv9Q9JYQ36oBAgqhDYiZ0N8W8y5S1d+hgp8X3YyBG0pxj8CigRkFPd5hjy2iymsIgfMAgd0gAUIgDE8ZizkQiC8wSSUgxfk5zHkIw14GkKc50J8AeLtwEQ+ARM8ATH+GT9sQxZsQ01awj5QZkTepCXs3xCIjTsQTb+h1iOEQGoqgvRggz8oxCeEAKyIqKHIg2zKZhbEZgZ0gp9RgmVa5k0yQSuUAe/5WRmmADBkQCxYQPQpRAdUQiU8wRtkQxw0UkiR/6ATRZXOJM3iHdMkLMNCOJ9aFsQigKVElOdnnKcxSUQ1AMAOnGPjMYRFsMFbcoAfqAAAAEAs2BVo/UPvyOgICEAkoAAChIICKEAC9GkCmIAJJMAhYAIAYAIm7MAOWIAKxMIFVEKjXkAuMEEJ8MIqQMCCNiTv/WQwWMLeLEQyeIlnqkR34cKIJtvFLcTFvcMP2ABCgIGQWNw/4EI4kKQifIIirAOsioRoOoQ8IIQ8tCiwtugR1CROTmYrGAIfUAEvyAOzZkAhtOiK7g2X+ozoaMAwzEEiVMIeXIAKWADi5VoP+IhCcMKmcWP2cakjham7PCL1kQTSdQSTSoSWLoQX/P9DJc0cQtAMJYpgDi5EQhENzj1TlErEIrCBZMyMH/QAAPijiUFjYMyAFQyljDQkL3ABNGjDnibAHCiAG7Rpm77BoVpAYRqUoxYpCxwCG+yDTd5kbm7qPsSKQmwDCfxDyzBMLoKEZDXExfnDI0zJAqwDR/7KFm6EsIyEs2ZBQSAt0spKQvzqETxtBhiAIZQMPxTC04rB0x6BGEDrs25D8xyNA+yWA4jC2JaCKJRCKLhBCZQAVTXPTKRiRv0D/NHMIcQVQvRra4VZ37GWcYJEdzpE0eFtpXEpge1AmD0EvkASPIqEWP7DOYKEJboiJryBx44AbxhAcwDDMAKHxELsCET/7AhM5Nrxxj60wD7wwj7Mwj6s7uryRhueHIyeiWsyGM/Wbhf+w6mSKuwN4IgCCtIewT9kLdZCLRWUijzwAzKIQfJiLT8cwSqIwxtELwD0ACeErfWObRfIgiyEgumyXSvkgiGsncpyQSKMABCwQAswRFgNChuYQrt2I0LQIOCJBM4pxOt4xuT9QwFAatweU5nmq0khhNTtQJsKQJuOwD7wA9441oo52qYQWWAEQyvAqCVQQgXzQl1lcKdgsAGg7vFuwxH86j/EJkIgbbvggqniwqmGxO0ixAq33oMA70K0QfEghBiEiSXkQg5TggevwnGwAKqMQBTkAiekAzQwA288/2ZEUhenMutMuF8bAhvArJk6oquErC8eDdhISEDsXBj9/kP9FkQjeIM3PAQWpwurqcDAmgtWKgSrjUSbKurubAMIgZDJMAQDy0MhIAMyFA8E/MMfF0QgA3IfZ8Zmroat5GxHtHAAIkTQckQySMQNF8QN03Aft8EkK4TyIoOlOmgK8EZwdoood0oHf/I+8E0h8I2DWsLUHu9MCGe8LgQmwi9s4C2KeJT74DI1uRoI4KuFFMRZFZFKMBkhzGtDRAoALA0L5MAUqIA4OGiYFMTsSsTMNsQg23Aht9Yu4q7R0TBDeDNDXLM397EY3PAkm3BBHEEWZO0R8IMYyMM78cLhcv9LQmDevPQtLQ+KcGWGzRRELMxz5tiZZ6BlSCxeDkiAFhCwABDCKsjwij2ErGQzHt1sPhONJSOEDMuw1WotRyPDEVhHFYSxQuCzQlhpRaugqomdADeEqyVNIxXE5MGfROCOi3zGHQRA0SDXUXiAB1xBHiDD/jEEOjvENfdJlITqSTcEONewShQ1QvyxN1vyEbRB1lL10z5rFbwrc4KESVvUSxOiMHuEvBrKAAydVbHWVzfEAP2DByCEB3BCKKzCFUwz8SRENS9EIN+1uTxyUusMBEBAG0AAMrTBYIsBJnOyiARNI+3CLvRyQSSScXpUWkvILPd1QZx1QdzAQlCA0fz/QxtbFAzikTErRD+HhPLICtM+NSDj9TeLxDqrSMaBBlKXi15vRG0LMglAQG7n9l8LtmCDAj/Ewg748lY/BCHsQtJ09Ums9aA0omWDBHHHrz97hs20HEKslUSUSF96xiD2iS4IVyNVwRAoZvFUqjWvdkEQNg0fgawMNUanM0dYYZRok0p05kN0Xf8VRNAiQWZIdEg4NUOQgIAPOIHrtm6DwiochYpM9nM/RCAETXSnmrtNOEIUSEPsgi98dlOtGUMwOEd4WUh803aXi4IXN0gAgoMVxBc8k6BECgo4BQJsgwKsQjoUxBzkAQSsQjYbdtI2xNY2hJDw94NQNJeIRNGK/8RSh0RtEzgJgMKAO7mT58GA5wEdxENnhEJD4LRKNNPfhoQvfEZGNrhEqNo/TINoMQQN/oMXI8SXOwRjMxJHEPRJjHj+ELcmLsQf/YMwd3mJS4RmNwS6BIAADLoA4MEXvMGgowAhEIA4EIAcODoBEMAZoAClCwAIYIEHVGo2o3ZBFEKvdnofzyIjsIMWvuq8wEJCrACiNYTYdMRKgnNv/7FuCzIg7/aTM7mAO7mASzmvg0KVW7lExLJCrHlIRLhnEIB/nkSbi/lC0MKFdXkZS0SaJ8SyPwRnL/cAscSJ7KOFKYSc/0MYFISIgPhCLDsNRg1An0tC1JoA1OUlYME25P/BFWD5P6wCKPh6bl8JBFyJDzvBDVBAJiRBBVRAM2ChMzSDFDTDP2DhOaxDNxzbPwg5oKw6QwyCQzi0Q9swQrQBCdABKFjHNsj1bq/Cbud4b5PAFdg6IzS5r9OBy+eBXBPAM7BEALz5QtB7QlQaQ9zvtCPEIF7CLjTThQmAh6tIW3dEAHy50lvUtXcEuqS4RLSxL9RRX1b7Q+D0hRF7Jv5D/tTRPpMEc7e5L2h9uWBBuI3FP4gDDqg9DhTCFYgAydv7KjgBBkj8Pyj8P5zDjP1DBeBYQ6wAbLgXPdCDHuhBM6wDPaC6Qyi+CMiKPADvJPM4QvBDeiMEKCBDMPgCY2//Ph7QAAqcQUGA/guAfkF0ZXd3mUJoeUik+z+oPkM0/T98edGrSLKPhIaLhHKHRB10Gkg8fX68TKapO0LEUUjcOUmQtEN0vT52BHOThPOV12KogkkkRLgrhCaO/T98/ll+PgW4Aq4mRDMkfkJYPKMMvkKcA0dgYXsNguIjBDU4wRVcwR4fgUdj8j/wQ5IrxEXPbBUARCABu1CcMWhQyRkUNAL4+vcQ4gcCEP8FgLiLYsaMLzR2hIgFg8ZLHil6IAmx1r+UJx/WYXly5MuHK1HKtHkTp8ZoDxt1hMMqYzFvOTOG+YeFqExaSZkyjcOzaS0a/xxe2qXkH9Z/hG64orbi/5yUTCtW1ICVJBMsajX+ndNTYV0Sshlh/YNVQ4+eZhl/QOxLdG8zPXIH/aPwDwViDFVuXMmzahUyyRCQQWhjGUJmCCQ0k6iMjAQoRmSqBAqU9d/UhxiQZiRHVNzLnhldZlTdFHdHHBBB5O441WFHjEk1sVwAUZrNNSfTrHmksVExiDpu+yZ6xqP0SFFpkhTy8PBElrogAspovqOOnGEouDKz5WEFKcJWuFr3rwLJ/Ofy/9vL8pyOnPlvQGf+MdBAAZFY4R8MDkPsH6OMysiGf3DAwYNCrtjGiW2uuAIyRhR47LFVPtwGBwKMimkM2loKrhbpmtpORqhYCg6nG4LKSP+rCW/SEaIa/1nKIRytY2k33I57KA2ZltPoKSYzipKi7h46YcgjtaSoSSpJSqmYlIycjiIGt/yHG41U8SgxIcgJ4QYR2HHCFTPz6+8mPE+S4kCI/vMPJ7LWEcaV4iCqDSIg/3HFMMPCwFKlIJeqZaTEEqNBCBqK/MedhwQhSTorb5Ium54aAcS8734rRsgjW/yUx5dg/afVmbZUNdItM2lqDTgg8hWOnTTy9cwt0UPnnzWZe2mpGquDqNOcvGQK2YdkdMcJEf5xgsEkkvAoQIj0hEgYm8JtC7cKknCFnodWwIAGRDTalST4KJJuKYgg7UheT/8pTgkldMiXolGSUgX/PZsI9she8Gw6AVecHtyyX4oQUY8pPoulqIF/nlxjGo86vmlhiHjYl6hdZ1Xzn2uywcmOk9ZcShVlI/jnl4waZqrJnNBJJY4QRHDCBic21mjcI/NLYpAa+vtWEFV00AEJiuglKeEhlaWFyNT+kVdeZf/BOCOxicq5YpxUW/PleikK6SGx2X6JbGb/QcfsZPP2KJWyvyx5XoogwfLPox8a+SZWWFkz571xIrjqhzZhSZW+DRc87Zeu8Y2VNIB6aAEn2PmnQkX+WeHqf1J/6L6kyi0XaXL/eX322mVKIpxuIEJik0yoYRTlJSHaWaNq/2kbEVVu/kXZyvV9SAcsNXac/yjLiTK+KeqZAhyizSlST4rIZbr5oQgQyZl7iOjlISf204DD1zUQv1wjbj5/ifyHeLhfeOE1gmRN1vvHtM7Utxjw7CHwe4mw4LCGUbDDBrb4xx8mCBHUoW5XutPItx4CO4ok7SWt64gwBvUSdZVFhB1klCtWZ5PNxSEVaUrFDDUSg8oRkG8PgQSfhIEED0ZMeznp25qqhY6cTU4m3rsJriL2kJxBAn8kIU9GUrE4jwSRfvR7RBp0IQ1ceFFYJsvYP6QARY2QZ4oDFCBEYvaQe0AkGsCCCA4hcgqcpPFXTvrHNxrQDSf8IQQZUYTRMsLBQoaDEb2wYOuQeJL7xMVbTf/x4EMMmZF16I5BgxiEKyBxP4/05ylpOuM/WME+/YnRLxAh3xo9sgCNUWR/pLTJDyyHx3+AIze4/Ef+MnIKXlIkcnZMFkvM+JC/nAQXGSkmD2zZFFw8AhfRbGMWNTI/Nu7xmqQU5kNKeZMICNOUUPpHcqQRs2k86SUhS+bnREmeaCLHH8L8QTiZ0gD5eWwN2DBDhSBiCwnm7h8afEkmwsGOfPRCkR35g5k2SMl1uYItORHhJCn0D0WSIh/JoMZYWHiKef4yI2j8HB5ZkRxSRoOd/+ABFOdJy4f0DWhqJMleNJbMmCVTlh45BS4Ux01pNPMhO7kZSDNi0pv84D/HHCX/RGoJEV2wzx//KOZLqRSNmJWUIqzgKf6a8QOizsg322lKz/5RBJZY5CRKpOY/fLUMLxDFJC+hUgEoIgPfKAAVG4PDNJlikmpQZBk4MUFOwkiRJchkAA/pwFpxspMSPCQHD3kAY18ysS1pQCOleIgKziRW+gFAADcJbVKwR1micMImBJQARBJDPyL4Bq2mJQk6KZLMw/5jCSz4h25ZIh7ZasQPOqAtRXhLkdlApB6/Zaxm/6GC3iiXKKMFAEmMSpKh/OO4aoVuFuMwXS0poCmZ8wge2FoRiIz2JHPoCGc7Utwj4VQjFrCJHyBC3ywyACII+IcfXjDcaSSGBY99iBaw/7td+mHWBzLhiIFlMomTtPYk5O3IcA1njY0tgiXc8G5H7Lrd2DL4JhT2yG1BDNyw/gNx1iyxb9qx4owct8FHg0PHOqZdF3ckrkn5AFPAeyb23vhIQADyQ7hgHRqHuFj6NVyLEzzkKZHkGGeKyYy752TrFMANLCFWRTbMEmgQZWQftnJGRDxmj0xAI896CVkh8g3DJYCy43hIi/+B2eZupCNovolnmcLntYbWwoYj8cZckMW3akQBCQAvePPqkUR8DyLLmV9kCewRP5sZ0//Q85aeY5NLZ5opib3cdrZ8Jo6Yda0w2BhqGdzoOTQaJ72yQxpo8QLdzmC3D/EFCuT7j//TBAIFKPAFDX4mKlDnZrDHvomQlS0TDD97wnRMq0Y+faY7aETMzd4unG9SCdb+4wWB2MEOqvFXjTj4IQ7u8j/eMIWMcOHLVl63tjOC3puIkiR0pXdGRP0QDGskuR1B95GOm22cREEjEr6cqsec5Zz0+CGwpojD/3GBx7J34BDJeE4OfehqlOMfPTAGZLOoYuaoOLFo7reZ500UAKAaxIU+0wD+zZLA/mMS5saaTEyelChf+9qXm+y+j0RXPpRgB1t6a5Tf2nGQn/sf7u7IE7Z0ZJYIQMxwWzmoFc4UVdi7IzInOkRqThHaemGyOs8JjMfukZi0XdGLDgVFEsEHzm7//ND/yLtvbv6Pp/9j6HqfhBcmMQUWtIIFh330mdQMEQB0XSNbB7U1yiyTQOOmsExh9UPYcCb8/rbnG7P6Py7/kpQoAyKRfQjF/7Faj4D9JGIHsQKgEYohxCLpJ9k7UfK++5P8Xe+AH8EFHpILqu9486DugnWKbOSmqIDZOQk9Syrh7Yy4QPZz9s3nGcz2YmX+JUNxxD/Gf5LG/wP2Z4L5kcC7ig0c4se4Yfo/oqyRv/Y+KYR/yA5YcIiH6Dv5mKIESmDQ2o4k3uC6GKu66EcUIELOkiL7KGu4Wq7Eyo8l6mat0KkAcWMVOOEDeu0lci7ngo8oQK4cRhD4bgLk/soE/0eArrggAiPwJspgCcpgzLiPKRJQuaavIyCM+F6iHVrsAFbs7UrM6p6i2joC9UgiyxjOJtYPIhglI+buJSCvKUzhH6BhAxIh/l5i9wQgtPruJe7vH6phBCni6TaOBM/trQBgCjoAtQIwKWzw2JovKYytKXqA5/4h4IiMAwwwJ46BAmVrfqLE4G4iy+zKCW/iEiqPCp1kTFiCgHKg0v5BHHrAC3xP9yDCCwAgAIpBAKar/mTiBB8iBQOrFCHi71IQ5ygCAAJBDjjBBbCw7ADRFrXNFGQwKdjs2JLQrKKvKYBAyJQhACovJ4bjJnTwIazgH1ogF3ZAE1+i7zBB3R5C//9Ywgyz0e86QhPFECIC66+8axIA4A4YYBHYoBZt4rAEzK5yb8gYYBb+wQ63i74+TxcNZwOODRNkQhmpCYciodSySMQe8RFxw/88YiikLtduohq8ABxVEd0aMhVxwhubYhIqEgCiwA86LykEDCIkwB1rAWRW7A9XTPKU6wENzBhZggePJg2y5iEsYiUz7dH0TSaAQAJiQbfK4QFYsSOOwSHpb+/+qu+mywwfQu1I0RpRMSjLIShtYhLGsQiI4A+V7HBw4xANzCrHDgdBDfzOpPS2CxBmMotCQb2aYvEg4iBPgup4L+e8wCfVLrRCyyLWzcEOza0ACyICL/BA7q0Cz63/ijLd/iEjYyMjRk8mJAAE8VC2Nu0hutLA0tHKFpGxIMwmLELajoQXh0wBIC4pFssmWADXXiLwHmIKRoCzNHGyonEEj5IbPWLgBjHdkhIMKyIAAsEq4QsrXYz7iky8SKILtUQybQILfSMfj0TiSAIIHAEYWUIPPe28spIotvIhyBLUyiwtPQLGTkPqShMNJQsiRsASVEAN/2EfTXAw/Q4uM8InubEcBBEAQAu0sC4A6jMSAiASiuE+oyM/T4Ui4sATcIATKGCbSAKLMA0SWpIi0m/fOHJLkjMnACEgMwIKyazAYvIWcwNCt6Q+2e0f3JEkbs4LVIAFguEfRiAp2VMV//1u8JpiskoTLpcO9arhGGiURjEhPtEPrSLBVPCAEPArnHqOlTL0TMzmsNbStEryH+4xJ/LKM5NiQikiOE8C6/YNSe8KJ0DwMtmtB0Yg6sBzGztCIUdgCh7AO19TI6LxJF4U8MBz6MwU8OC0J3vS78RwugBgB+TAJoZUJiCTKIinKRQUNwQ1KfxUIwTMJv/BQeMNJ77g+lAhrza0KewgMYKOJTaTSIcsAASgS0HUI+a0HLwUGEZuDdV0Yx4gsCrSFPeyTUkCANyAEIpJQe2KCbLIATIVEGFNUl8iSjuiOaWEz2ASV8UyAHYgFqZAIW2CF2KhI/rOVH1jssqhHNwNPf8/dS+HLilV4Bm+ali79UiQFAQYtMeeFMweAjsewvU8QsQSxjr3MNMK8vusQQBGgAXac1UhQhmYNRcAy15JIkVZojSldQpG0yOWMCPgVCPiMxByBjfewHDgoVAZzL2szM5yYu7g9SSYTSFDpiMo80zWsi3p56+Wk97OdRrSAARYgLOU4UzF1BAMIepadhU14kx9UhmWYehSVe+Gbgf4oCNAbgrKQQ2CFid2IX1kQgX28STwy1BBrFYNSyOSJENbjM6a9CHIlSIq9HIyMyNeK2SjCyfQju5AbbGmKBuiwEtxYgQ6wWelNSdMsEr3zguQlU1b9iFO4x+CYQTKwWBR7zT/DSEWvBTkUM8nvUsAjpYkOkz1honfIMIxvbXTvPUfuC0nQPArIYL1POZIHu3RvpYkejUnUHXf+uYbLuEZ1ID8UpcklAH1bi1MiUIZqgETRvEBpqAV2pYidgB17/Uf0KB3OwHXDNZt0cAQgiEYiJZ3OwIAfKHUVIwbFuwhBCyyHHZvHpeyOEBJbeIHNxBXh7BqqelXbUJB2xXUnsJuPYJyX8L1liBR9ws05WUNaKAHks4CM4JwIWJgO4FMWQL1hBdhEfYf1IAPLGEN23QGvHTopsBE89YSDKFM/wEI3O00H4IKeIEKRmB3VRQpKQJ0M6LDiNThnvZo5HCttIF+MJYl/xqhg6tJj87EpCqPa3PjuXIifScMXbkXIgghgQKhB4RssirxZx+CDxw4BfuWVYV2BAI2VAl2WiXrb9N2Wo3Xd4k3BWYg93x2B3DNEHzXAKpAbxtsutCBfD3SFic2i5h0zF4tNwASEL2PIvrxcpbvIZKNJDhWAg6vEmSABfAgG67hGgBhTcgDKEYgfEnCS0dz6HwyWrOYD6C4HLL4H6jgRE0R5HbgNBp5F6K4FSAiGIKAF3LhNFvBEEYgENLWEKggA4ABDdDARM8X56LyDUrrJUQYJ/SMMaHrB0mCub73JtBYJkBTJnIZN3asI84SIrBWCdEvqDjUjXNDT7UMN4DZOv9e4R8gNilGIBcoQRx4wQ9iowpQIA0WwBOmNCOAcQQa+R/6V7Kejk6F7yFGIOncjZWBQRxKw92WcApiIRgMIRB2YRf22XcfogqAIQu8+CFWeQZMdJWpQBL+QRIMgJWlbvySFSKPZ8vI18qK00LnRwaIb1+pCZlJQpi7jSnSJIZzYnEv9CSu9CWScPUMTBmAwOGkebt0ixJm4MdGIAdYYASY9UO/tJBNM/VwDfiW8AGwGRP/Nm8fYgZ8Fxj+oQqeoTRMcWBN1HjT9qAXegiAoYurICOmmAqGoAlu4Q+G4GWRFX+lbnBZVAVUoJ83xR1owJY4C22tY4ZJggAw0Nmyl4X/hYkJLuAJ9kByHfAlXuslJsK3XqLXwpIlaKAl3fik6acn0CrLiICmcQJTfYMSzDgjpC6ozZlg/a52a9cYqmBfAwFmKQINwloSmuA1oJpaR2CBt3iKszqsq+AWHBqqNWK1C4ERHkIRhqAKRvlDR0CUQ/tFa/fpqiHpki4QdInxQEBLTatjWAHhaPkkqMEWhxAffEO7mWKFNVO5nqQnPIuzfys4BIwXFvJLO0INUFchA6/8hEwNDjid8ddLn2GsFRoiqAAYWvsPyAAM/uEKyCAYduCcOwEiYBZmJXmgkQEMgrsQgMGrv5qhJeEW+uAfQuAWJAEYHPhvO4EXQnsv4fnp/xTSeML7JEoSARRlrTiAOiHCk4irI5hrsG9cIBeUQVeMvj5Zgts7g0dgNDM4dcfvRQc2bf3WRDP8IVKbCgxAElpbEcigEAQcDCY8b1NbI4IhrMU6w2+hCTzcwoeADG4htwOpD26BDD58BBbaAKiAoqMun7EaIhh2u0pBjnNiOD1ipHF8u9gYoxfUyhCHz/bRI7PzJNJ1Y8i4yPjAU4W6BLzU3VTgvdm0/E6TjEv7H9I8kqEcwzNcwzd909N8qx0cIhYaGIagtSmiD0LgoSGiCtAg1Rs6t0VdwwOhCZ46klE5CNDAS8vvnM+ZCnx2gdsOB/f8JvLgH1LyIYbh2Ez4SP+MOTdUXF01ThIdFbqaOSkkIAcevVjo6xDofHdJ1GeHtr5nwN2izxHQOhdGrsJzO8zH+hYCSSNCIATCfAhuoQqqgAoGWhxUnQpqPbc1vA+aYKuhmgq6vKEpIpA2IQZ4ABxyPdYNIAWeWsujTpR9V5Lzdqo7ogj1nK+BTLD9HDfo2JoD1Snc1ToigABYOicEANU++B8Su8TWOxFYYAp21xE4SxxOI4Jn4OKFTMjy2RjMvNYfAgoeIh8ogoIggoKiHOqrYKwzItRHvQ8CnMIdegj+YOr/oQkeog9a5Dhi4Bdy3b8zYOMvvr8TXtarABmv0iag+zH/4d9CPiMacLBNoIb/WXi7ntm0ECUpZHPMiMCwV0zP0OyTMZgixmAEJH0GcoFgCYzAjrromyLpRR3sR70b+mDz3aEPRmEMFoDDm4AM4gHpSSIZHsIJxkAcYiMLUqDCNz6LT5kKUiAI/iEXxC0Q4gAxzQsiSAzbScLuceKV+jQegawL8vwfQrpYHLTEGLtYRsYKHwIGpvskuBU3Mjc3rFn5k2ICZoEXRjyAhzYQpoAPyGAMAiHL1GBtO+F4/4HAmI39W+QhumHAcWIBRmEUumH/AWLMqDGbFiyIEQOcLju60tgBp+ifxIkTSVCUqAgKGDJNmvwzIBGNoRESO1H6Jy7IiBGBVgb7FygQpH8N/y7azPFv1z9dFxdJ5PAPqM2JGoYaPYqUC9KlTJtSdOA06j84kf4BMFpJalMT/15p/Rp12b9JQ2s2LSEUrNQAaqN2+fe27b9ZvA7NMDYj1gxDhnJR/NWkSst/najMCDRlopYpI4yhi2FQE1g7U+3AsYN5px1Wulht/ofrokWk/mz0idHn1j9JkiQGQTMiWCeJIININPQPdzBxY+ROZIDUgu+jSocbP96UrUQJUQ/IfRsXuXSmMIRPP1r14pLrXKNHzeVH6SyJs5hxISNuyERx/45U+VVlyAhDVCS+/JcYv7JYKHgu/EeZTVUMBYdErFyU2UShXcSDVGMsMMoCY4gjyf+AaFBx4T9B2AYMRRemkIsva9zjGyf/mEgRBRQVwcJFziEH3HUyyuWNU9pMNM5E7czI43Qq9Dhjdr69MFEZNhXH2y+EtKTGCDMAsw1MrHUoERXBkISfGlMEEsUvEgXYIICTTWTHgv8cKBEPAV6Ux1G68KDLAuIAg4ZNHabwDxVUGJBCBoZMsUMU6NhUC1g+SXToUEXt6MM/L/oWI5BNJWCTd01lZZSQS7kgUVGOGlWApNMtQ9ZX1kmqnHFYGlfCRH5JFOlEiBijQg6J8WFJLoX804Qk6k1U2EWMkeOlM73ZZKZ0yTKFmS7uTIRhfXlm8A+eGaRgABpBjOQIS9/8s0b/uEZp0RQHbKS14j83UuRpW1zEOoGoTeUIF3Jp2NQqE/9gelEpTB0iUbzyyvVAW2oMjHBTUUSFDhZYjtBKhx2y80drIEmUAnsSqaGlMc/84wtSaCY8kS66gNMEMNJq+NE/GQRRW55UBKHnCFsGsoZZ/xRzEbn5DbUIUBwkOpWiO+4IKawkIyXKP01DtXTUE/2Ix3UFf+XGqXJZI2mrrdpEjUSUSjfARHGQ0wN+89k2USHstIYnxii9xHEgz6gmNVMK/SIJlbZRkUIWeVI0s54zz9CxKhSpUsRXKCK1LlG+jRfUeMVJ17RUjT7FI5b68uhv3hQBIbpcRJYe6lFwnGHM/8HBUEHlP7FDcMVqtq/2zEtTTBHMx00tC+QCcP7yTGtVGpCFAXratCHNVBgSzBQWBALORKooU3pTlw+s83DdN9VIujx6lX3pZUt0jU3TfAVC+RMJrAQcgcRiMx9BqHwR2y7vatPHHo9RvTUxi0xkGplcGrQQd8zpI33CX5UosqHC6WkkN1uDRNDROIk4onTfc59vOriU8E0kg0dBBXKg5kGSYSB9NJmIBbXyBfcBBwESiZ8OYmGf+7nGTrIzwBA88o8YBOgXC3DHL4BnlDXxRCJLPE5o7LCAf1TBWn7TkP7Y1rzCBWEGgOqSBVORQStsMHtmaYA0CgSkR80IhEgRYf9UQvcc6bAxhVpx4z9SdZQY0nEivogFH/6BK9qsTHaDnEjcyBSaAyHxK7goExpDs0jQKAg0cIiBO8ggjx1eZJAbyhPNPgmbHaihS/9IhQYnMsY99mgYx3GACJACCU8ATCKJ+EcHJjLHGaVjIpnr0fmaQjpVLs1SYKHhRfiwhGDob0/G4YyBtLJIO4TpKGHqjMmiaLyL/Y02WLQNzGC3IejtbgpKAActlvJCYXqwXUshBMlI+I87VM0ooiDmcCIlhxYuBSdaUZw622LPi9DAKfGCQy3u4JdA6jBPypNLIyOJFOCVaSIGpChFPtMb9VxMk4OzIstm9k2a/Wl3PUBBLX7/9A9+jpEt6bzI4/5JMlG8sqUX8cRFZqnPpjxhOv6CGgpVCQOjaI0pv1RaVAQggIlg4h/wXAoTZDCRSxgFjkbRmQ6iEgaQITQ2lmCZRGJnE2mBtUfhkAs7tNLQj4B0Q5a40hSaFIh/LMEKMEUOVZGDNLB8QFRikcjpLtIFUfQUOQIDC3PuZRMUHKWpNoGKmYr6j8JqZalSMZJ0rqo9LIAsCrkYQSAnos0d4q+QA5vmUpIlsYtslCIg6VBt9qRFQ3DxrbFoFT+dYgqJ5LauE5GAMXmbsF7KaHtGSVtvkRJUiUA1VDLQ41F+apPffgUT2JMIY48C1aXclSI1IZFN7gAr/w6I9x8MUEoc/gGCXPBhBrbp6swsobJOAjd/Hf2K8gwQ0iC0Ypwz4AMfSrAdCdD1KkcJ2j9MwQabDFWV7EQOvVRZ3QX/A2rCTRh4sTaR5DLFlDah3FfYct2mWHZ9vmHB53aKlDjQwALqZUEn8EsnKljiNVXwZn1dM9rBHdIoofGPRHCxRCAjZ5tOuSIwYHa/PW3IZrsrwR5mgJz22aTBviEaU1A8kc1dR40yum1bjhHMoVR4vgnzQqkkVYoHXzm7xJEIDUAQi1zsxQC8qI8hOtRViVgCvxSRmLRAYryInglAninZM0uH30Qj2QCtGAHH1NCKz/2DrlLxw0RqoVh5Cf+hKbHQMJk/zaqJfI0pbhBdUmW03aWwmSJCAUqkQtYDQviRF/+AjSG6iueJ4Fp2vJ7IkWkjsh9b9EDETiLCFK3oGQfj0SVohVxTOpao5BNAAzVKUbQsl91G5QKlq0f2rlJdecUoRpL9CmLVAl0gAeHUX+lCqsHCiVhdBASByIVsLdHW+aT2q8C4xSiEsAkkCHwTo9jCFihAgRuIQ2M2MQMBv9SUJv6jG/JatMU7weQctOLJUN7OUuQtJlElmOEuvMiruA3qvI1ZLdIVHTwmEoHpXJfAYIHuyo1jAWPI2RKdQFwr8txrcWjiEWh8hAW/8QhvV4Ae9KgBBlzhCidMBIj/YKmeqPTnGmQjeYu7a9ITPL6Uck8Ejf/AqYxM8VJc/uMUKY8Kpa/jgHcnTSo7/aNNzo0ws+jEODy7u0S24LR/qHlGIFCBnA0xGzW85GIXEwcGfoD0iTziHUbRgyZsIBG82UI1IfiKGW5ggxuQYfQkNw7QuwqzPVvcABh/9AX+2KKlEFci3/qHhKXDiQS3XWrs5tpQ4p5uuQhNKih9waCEeYzehvgiNGXOUai8abVAViJ40PkMSGKFGazMtbyoghCi8QgSS8UWF+m8URxOkRXoYf3s1wM9AO8KHhnAAMCYP/3tH4Rlc2wGuUDx8pliAQQgKdNnIGfwBJI2Ebd3HIPH/yNe5hts1yMghxTVhoBSUWo8cgITEXtGEWZHwUIXwWEkgwKB4AZ29w/adzsfQX9NcAr2gAvNMBR6wBTmhxz0cAMzYn85aAB7Bgyd8Ggq0AqUUAIlsAMpdyBYdhGR4xtU5huW9g++JyM1MhwV+HFqIWnHVxP+tEcbKB0awIRNsQf/kGBWloA/YgGxcBJyNQOzUS2uZQDisAWn4A8wyBSUNxRUR3VtgQE4cB22oYP3N3/4dn0cswSvglKfxgoGmF1hyFsL0yNXkXxSUYTGhRRFiBQSSBEZyAQopy9S5RRIKDUdaBQfiBRf6CMwYXh/tARrOH+g9YajYIdN8QhagTdDUf8BRkEPPfKHfwgbTaIGT/B6EgEIQ3FLRuElRsFlUpEoG9AUZ5ByNjUjx1AqxxCJTZEY4XYRq2aJ04GNeycpZCcVztcUSfUA5JI3LwACFrADxhALLeJZLaMxKdAEmnCL/5CLuSgMknERs8gjFSCDsKBwxxE7blh/81eQ97dFamAFajADF+Bs/zCMSME1pAgkzKhtRwGK5ZNLDmYUkyCN1dgU6igRDzkjNPUPTwBVe4cHbyBMFygRhzgU53VKefMjKmABcMYHVuBZG4Unb9gNMjgICPMt62ATZaWLf4gt9scLhuCLqwKRTpGBQKJ7EjGVIucbcSANkoJCNycRIMkUO0D/WRPBiDbxBtuoFaf2BMCYLldBc5KCd0cxahQBdsehAcnod//AhUyhAi9gATc5grGwijMAEimAJxDACEcxE/9Qj/8gfv/AAxB4FJ1Xi0NRexUwTUUUaL4ROyBhkLtYf7ygEo4GMZ3ljRThhAnDBo9TlT3Cj2k3XeWTfF4pFSgnERlpHGppE5jAkruXU01hii3UAMHJCoHQInOJFC+wlxbAl7tQbyfIB9uwChcRA1FRexYlFRQ3FPzIIDg4f9jinXwyf+JgCYMIMZSQA7sQByAUL2InKZwihr6BbUghgLxJEcmnRya5FBfAbWPpadPBbVAVliSDnzYBkzZhFgPKFBqA/zTCdQ/BGZypEAXMEZdLkZw2iQK7YAziUAhG2RbeJRExxyMhyAMNYlpqwZlJCZ7f2Z2NppNB2CIyaRMtkDerGRXMqAASETZN4Z6iMwVv92W+QZvywma7+WlsJJtTJjkX0aAOCqFcuGpGsZd7CQK70ARSF3MRAKJycQrCYGgyMk0N4g9p4hspSqbfmQKUMAMtygtO+Q+JOREdMAHFiJozgg5pIJNscZpywZJEKjV9NRFRCSSmsAiuORTOFoa0aZYXwZ706RQ5kzMNoAo9YJx7UFgGBhRRgJw3GRNOUFZe4qnSEQIqojde+hVmWqYpagmx0CR8kAiUSBEtMAC3BKcd4P8HnsATa3B8MjKVZGgcYelcfsAGNHoRefWbcpEfPvoVyuCnYHEBtnkUaYEuGLkv03oUF7io83VmTCFcjhqckVoCZeBxTzoRQsGXfGkM2xAOXjKdFLGuCJOlw9EgAiQVp2qqdHYlEMMLLXJuEUAEsOoHcRqnlsYNNiF3csEGLkCox4GNF+ECzDgUR9MjloisUdE44YZHTiGuWjF7TEGFEgFeDICJdZWtTiFcwfmoiOAJJbCJ3PY1kmVg/1CuFvAr1RZETdGuS6GPyLEJomKmhEmvwHCvrZCvmUYREzABLWC0cSoR0UATShAF7VOwYMEGGzC1PlF6MvIqpfgPSJNX/+T/XDziBqnzD7XUFEEKSBcBkyE7HCEWKmLrFBupFYnpoMGJCCxgJLzQAhfAArEgWQxwKJ6AnIFAiVLwoRMRpuyKFPo4i7igndPxAzzLJz5LmJNLuQYwEiOQCy3AhQ0QAXIwAEmLtHDqCXDwC1jAAiyQqNLhnjvaFl0bFS4ZNRMLXP9nE6FidwEqKsqwA9iDu//QfwPDSmUxtzQAA2VACbyAK7yQXZQDshwwAYA7PXfgBBgwFDcrEdZbs/v4D7PYuKdQons0mNXinZRLvimwlE7yD7zQKnAQnPXQuVzABUhrtJb2AYTQdbHwI5njukvDbVVpl0aRp6VjnG1ZVwF8FLb7/zMXsbHIwbv/kLpuKzVz2wAnEAtMkAi09g/OxgXxohQMABQDAL0xwT+Ee6UU4QxaQXmUx7gSccJkVr4pMASTG8OEuUUzQAmaCwJp4KDOIAfwOwEbfLSJoAI7UA67EwuuWj788g/Fukepqxa0e3YHtm3/wG0mCCSxcgcELCla7IEFUg8N4Kg04AYlcLwUwQuUMx4gOwF3wJcxESWb8K5fgZ1HwaXXS6Ix8L3uA8MvPMM+W8OUkAgwkMMmKwXhscF04cBT4AiKrMgzUALFoaASEZ9tUVFOIaMyMnhMrBZOfB286humwLpgeAFhyAcJLCoGrBXXihzSEAfgsAbRAAgq5v8GTHC8aSgRNswF+/AuDLDGfGl4QxAlUQQkYJomh0tNjikVjTscMXwtzbzHzrxFycsCg9wAcKADA/AuyKsCWqIGi+wI3ZwX2xAPErG/QIILjui7QOK6kwwW7DZCEuGAUSGK0SUjnLBboYwUY1nKdTUAuwUcBOgbwUsRAeALeIAHL3CAF8ALtPZHX+NZucAFszALd2ABU2AJyPsr/xBFXhJz69rCxxEmI2oTjwsJIm0UJWrMsWgU2DsU1OLML90nMb1FQksJMoACjxoDzyAOf8QYCskxb+XNeQEcGlAKjVLObYGJcPsP7NwWD6YBPqDJSBFMScVuULwUGfR/MTIAanv/EXFVLlIBwRdBJAUqOgl2Lrwcp24gAAEQCY0wjI2QHWQxslJRlphgASPgkHvAC9rQVnI5A38NSBdwwbPgX7HADxRBuCtduGrB0hOxAN3QByFAdYoABhEhEWBACmcFBhdB2cjh0jH90kOQARkAEkJrCRfgBjqXC/Rzyyuhk4/GzVMQzg4gCqJQFFGNc0cB1c5x1Eixo8F3HKQjAF+LMASoKRSBxAgDspMiEVwhKUHjvHFaAEmVHRHpzkjRBfZEWRagDBbAAg75BJSgDXz9Dzh0glAmESXAAsfbCjPQCrhSOxJBwkbhDI1tHJj9CRMREfm93xdhBKQAJC4t2qA92qQd/wy3Rgn+dYL/UAZ/zQIzsAQj8NqP9lZTwAd3gABQc9tZthSVTNdMcQBP7TgTAdy5fWrXDSRlI1lKIBHHDSRjuRRC4clMQbbD4ariBbIDUAB4wNaN4NbtRhHStVRAoALf3QrNygWrwA9DMJ56seAScbz+xQftTQm1MwoT0dgfPSNGkN8XAeD/8OUTYQT/MOYzQi0uM+AFXuApYAhByIYTsV7r9ddpCuGiOQM8Zwhe3SkUwYBZCS7/IFVQ+BWNo2G0OQxF4RxaxtUT0bD4zC5OkdxDQWAoLhdFIGE+wcuR4owXMc9OEW9KlTfkQwS4twiCagrlNQGJgAkCwCVtDdcC4P8FXvAPsj4JbEEDN2hCNjE2E1GW3c0CuaCfF0AJSZ5JKTCeE2HDCe7e7t0J1NImolLmRvEJ024Um53fpNALpNDl10Et6kEtfaLmal4flNBV69Xgcj7nc+4kP7dnVJALElZhqaMLDfAN6PAGLPkF84Qcjq4V/J6kn4gUABBDxB2B/3AokvWW5qgVF4kUo5zOx+HcEU9LyEEEnHAoQcPLHVAEGJoLnRALuxAAsD4JsW5mARA+chAK/6AAc7AUmLADO1DkwF4JF5AL4n3YWbAN5hsMwRDlfFAGVJ4CUbI0O3sR2GAHMYANYxARlL0J2EAR+60I2GD00pEFZ04RVT/aVa//9ZbQCp3AC++97OvV3uulF69zLUnJC7kAAgnbNHPgBxdQCTCAB3bad9ZB8E3BknmJMAGF3Edxmm/AxXLR6TYxAYveI/rprNIBMAAtEdUA6RMhqIugxrygDKzeWU6y2lMw8rE+CQLQCChQNrmeAAng3BLh8g78BS+fUrU1hHzAAo+8ChmwDaKdAfuApv01A7LRJ/8gOMO8vdkJGov7CNhgA5b9B1LvoU/fG++g0r7R7RKRBb+i9RmA9RlgCXzAC5TQ3u+9/VOevNfCBTAsCTBsDGaZarxQAJXABCqAB74AAIlqyhdR4xTBkuYtHVSLMHw6HYM/FACh5N+/SP8CDBwI/wDhvzcgQCyEuAjiRIoVLV4caALjRo4D2QzkwGGWnx0AAOTKNWPJwBmtWo1QJiBAJBQDQqFSoCBBAhM85xABUK3aG0w7dqgosefC0gtP+Izgsopflm37LM3AitUQrwwQQf3r1rHjI1z/3plFeHbiWWzdwAxU1Ofbo3sD1/17O5BdEnuPxG4csjALwiyFM2Q5/C9FJ0OWKPExxKcVZEopDl/OYDmFvFxv/nGaWGqcqGFzOlzI9STHFwv/Wg80CtGUR4SvPQ9U9lf37oq3abvgHVz4Rs87Ng4Qe2H48n+T/mEiyjskAz9TAAgIdIjPjBFqFvJ50gP7kFDQcibQyVPBIf+TQavtUIY09dICTVkkisqPWa5YM5hgbcWyf7paCBQnFnKGOWz+KWugsho06xuEHtlkoT+c8WuhH/D6x5YEmfurMMQK+4cXQ7aipBMqDOBFHsNcHDEDGTMY4Z8i/nlloFL+EcUBUUiDJhHUWskBEwsw+WeEQ2KZ4h/juFiIDRcWAQ3EgcqxEqPbouCFNt6WYCHLgRAQywsvOpJooQnEesLKHHdTaCAkxWJDIomoewGASSZhgZftRuiuO++S5OOQfZgJhZOczlMgl0lMEsoopJSqjykWiOBCGy46cSmrTriCiMSBbEBogX8+1A2Xdx5hFcKKsHlkVWdCsIHUbiRka6D/R35YYEOI1BKLnY7kQYjYEbM4Qp4MTsxgqm2QlSfZZAsxLINtqhgIBNC6cKAUH78VJZRcmCCXhTd2iIWXXJZsEiEO/pnt3dkogk9MexfyYyHggltJTDJ1E+CfL+xt5R/lEHqoo1go6oIj5BZ6o5rgQppAhWpMEuADSoxBwxBA1QDZCpDVEJkPSriYJZRV5tjGGAEgfa8aC1iY74mmnhKHC15a2cOl7QIUcKLB7l3QVYtWXfWRBv6x458MByr6nwUpKouVe4WGVp4UqDAkBTH+kUeMI8Q+omzD+OFlh5ct4OQVB7j1sYseReGkUj74yMVPPi7gpcYdXgMJtCpdu3qi/8GH28G3f97laM6JSgjuRoruRODfjeK09+CFjEsYo3cXvrdNsaaboAdM2gMgFktyScEAYDoJ5mNBSR65O7wt4SV3XhIZqMt/WtgHeOBzz4WSVjiNzBLLZCwcxLL8mnohVRHyR2rrGSx8aISOGAhaMZS1pJNO5OGHn7HFML/sI/jZJpDrAFAhFG7nn9tHTopvgRfjJ8sbJV5UaN5uJHK4vyRuN4DrHIiAIAHJUQQBDAggRIzzHXrpJhaiE45zBiIx6UBQYO05BgC2YoAU/MMAQzCAARjDnSkESg0jsAJ37vaEVlDChjfUn2P0p78UpagTfKDCZgY0kMBEcDd+QSJEnv+Xln/4AxfRC6D2/sG97alPDFlIASUM0YkMMMN8ZNsG+54BgJLADxom6MIr0hiPV7wiAXPgQAsuYAiD/SMyvNgHF1DSLiNyJE3/+GMfBwK45fTgHwAcSEEQ4kHL/YMGG1Hkbgw4kC8kEINO+kcCN3LJ4ShEcX5kQCj/0YMdXOxlJskFPyqSwhSiIXbcARSAanhDHeKOEjuk5S0JRKyBEKgiXWHE1cjCoKdNCHt+UcswMQJFMUlxILxcCDL+IQaxDYFrVOiEJZpVPgggIxBGKSUARhCKNs4BFNBgBi9aMJlYnKhEi/nUPlByiFxEZCEMYIYgB+LBfemzcX/BA0Y8eBH/hWgwS4orAEI4GUE3/MMNLwAR48xVDUy87GXVyAUz9jERA0CkoyYMAhXQwJgg5MIxlkAp7lKauwyQjx/I+NpCihiqAJ4CIbh4BKyOyBFX2MtFA6GiRaSJkBRYwhAoyUU2cUc8lDhGZ48JBlZGMIPGdClsGTAqSpOat1hw0J8LiUK+BvpVjEAOIQETjhwQUrmOYG4haF1Omw7Gh692YKGOgwgTDAdICTLkH+8rwsz2gZiLlFCmAykfMhSrSn5A4B+O7eY/hvqPNhRraL6kCDTttcQliqWYurrpP8IxEFSBCFkYkWZl2/C19YFvdZTIBTZ7eLxWRKYVwTDELUGFkJb+/4MxBtjHzqhgiR54FSLvIhMhybrc4RziHzD4R5iUOxxANGIjlpsgRS44EOXwwQKfNOLAOCKDigQyIRv86w4kMAUV8EIMhi3hTClSQgJNdiCOvUhlwcZcJTYxONVDSPSYKaZoIeRr0pysaikrTVUiAwLl28Y2XNTSGe1jRoP5aaj2sZjNiCEDJlLXcvE6EC5AiazZvYhZ4bqcAYy1cCieCOiEw4UPbORNIIrCPSuSwLWxIAc5UEYuMowRXxbiCIrliH4HElP+/vciTbPDAhQhHFPt5gj6RTBChqpgLg+ksmObZvcI+4+hUeUw0VpfBoCRtxoZ9yLgLRwDGKfPh2hyIf9mbbJuPoBiz9xmCjAoGEJkzBwH/KNhDftHB6w03Yl8EoA/BsIUdiCObcxUvhdhcjQRAllN51k4AK7IlDdS2qvZFyJKVvJkxbBawhDLRc86ArTKxo8Pq+tcYoEziMTxjzV9dZL+xIFYVowQQHDkA3AemJ05YmKE1FiQ0O2IZ3Zx539IQAVTCCEKuLCN5VxhIvhdSKavFoHgrMCI5C4cMtqg7omgGiEKpqyWw7wQaY3NiikYQi5ssxAEMHsgxuizpwUuJhw8rCNpgFNF7jAQ8naEC42cSAIggmiB9+sfQLiOMbaxikoXMTCYFQxFvD0QU8ubzAOPQQDdIUhwU6Tlm17/iH6vbLYpxlp99i4Evt0XJ2UPfCCFXsgruC0mFPh8Io1AOMItMgB/L0S8E3nCQjFicIyk0ecSqDYlA4YAD1yB47t5eUXCbnSyhxsjbYB3vDsyWXZPExlHvrkVt5GBIRhSNwp5+tPLrpueG/EGAYyFZzAXsIDehq66oTqIImlEFaigNVv/TNdZRneMBPW+Cxn7P1Q5xV4yN+V7X7u9TA33t4uNbPIYws4pkviJTDugoIc9Rf5+kWEnnCODFkvThXOQ3bAeIQrZxRtej5AcLMTZCOm6Aq6w+fxaBNzuLtwJEILu5X5+N0LgLwku72B1q/vI6DsCxwG44lwPBDlviFP5/2N/kYT1PYKznwhaec8b9FPEM9C2l8T/chD+L2dgT8cDxSm+6/KAf7iCS+s0iMg8o0sQ6sszJNCNkhsO7YOACuS+dXs7mDoCCNiGaYMI4fuHHNOSAKy99bsID9Snv1MrtRoIQoCIFZs/peuI4DNBRZq/ioCoisiF4/vAf4iFMBELD6gCX9gFCoCIobMSZ7KSCKiQiqiyq5ECUgsgJRsOCCABCFiFK6jAbsJAfiABcQiEgeC9gNoFAdC7inAr2CtBi1A/ikBBjnAu4VjDjnDBM6wIINSNXVsI/NsN61oOP2DBvxJEhFg4jIC4itiGI8iAQiC5i+A0tSM5ywuOCqiIGP8Yg79wwI54wn/IxK+qQJezCAq8QhK4givcQgfzwlXAFsCRP1/oiDkcCEWziDMQJDx4Q44ouoHIxeUgAoE7AwF4Q1gEEW0IOo5YvOEIxIV4PT4MjjiwLhDIBS5gLCRzvseCCGmyPJCjN93YRIwIgVH4h5STwo3oRBARt5gTC8fSvoHQvnYkgXd8RyvUwgrUQlDYhh4IQyPSPxNciFvkR4qwu69ywYogoCZzP4oINoootrMKBGPYtjlYBRJwMCukSGsEN+9TH1GhCEmkiCeUPuZowpQrR07UxL/gHn6gwr94xH9oR5b8h4iER3iESVJcBVB4BXEQwYF4vRtcLn9cLjv/nAhoK0Se9Cc4mIhHuohLwIgeCEjFQcoAykU/HA49VDjmiIOFTIgiAAELMI5dIIRtUIBVoANQAIWIxMIthAC0E4O3C5F1XAgIFJNu5AgpEJOUfDeOcMuWjMm93MtVyIM8iAcFqAiiHAhPAJg8i8N/tBKj/AtfCAA8CJiDgKuAHAinFA4RuJqnFA7K/Is48EyIwAQjGRgBeAgiEAc5EIchQIAruIJQuIKyXIXYlKzZBCr1yayTgwi59DkIvMSOSAaxcEt2vDy+JE5QgEfjpAM2ugig/Ael7EXFhM6L4MGLYEzecMWFuM5/MMxCLDqldCSfJLrl4kyxuMoAEIDzNIki//gCPAgAFCAEAiAAcSAAOYjPKogCPEABFAgEFHgGCrDCUdxCU2QyYmHEfygEOjCDf4BAuLwaWAARG6DKi8iDatSvltw04sTQvcyD5KSDPBDMf8DMwXxBjsjOfhST54xO5pjO3biE4Yu/f3BRhAjD8dRJe0k8N8CCGEUI8MrPf5g2DMCI6wRGsUjIjTDP8xQAyJQJ/oRPIojP+cyFZ9iFXfCFZwCGLBw5A+U2JERCMsABMiADCliBJgjR3RhHi6iBjnDQgUjThShQsSOBCZWsdVu3boIs7rNTZDBFioTH/4xJ45TJPACFPFiZD31FMTSIjvAFW7yEEr2aZEzRSBXIi/+QyorYBc0MjnyciBvwvX+IgxG1KAGIBDzAAviMzyEQBxwYggiLzVWwSAa7AhzAAQjFgBDIBE2oAClohgpoBmeQggpwhtEKC94IAX1SQi/bNDqgg3gkxW5ChpfSQgeLVggoxVLkUw0FBWWlgyu4FnKY0oUIBRykiP6DiMRciO50PWHMknBtTIwAT0mVQYuIhGOsUYhCpIFwRUytCALgDSME0kSCiErdCCOczhv0hTfQ1IGgRRAx2DMYArH8h7LUvizMU2cdiCoQhgrg1WYYiF6FiA/Rg2H9h95UUEFa04vwtkLQLIg4sDbwQlCQhF0IhECogioYgiHg1tgsy52tSbL/7Fk6mANC5bhtEIe/A4FvdcVdwJZ/CFd2hYicZDR65deFyEHIDChHLZwCdNqK0NGKWNp//NSNoAWMEFiKeIGEPQjvFI4CpIiptYiyXYiD6Np/swhNvde/QDi4nQhCoAACQACwTACglVgt5IflQ4Zw0ISOPQeKoMQKSAJzG4gyHQgGFYuTZVOIqIE2XQjNnQgHdQKVNdAlm4ivyTQS2IZnAEZbBEa4CsMco8Uw3AUUEICFHQgjNMJ/OIMAUNt3hSSKIFgedEGrjU7e5YiEBZEiDaBH+kyLQAFNIl7dYFuLMMxIqi697QjDLDtCCASZDQRyIARxSM1tKAQyuIEkqIgE/3GGCqgBy03Qf5gyJ2AHM2jfjuBcNqWHuzgHjvUVPdCDf6hfiPAAD6CWsiGbeaNNKmyDIyjLKgiAKd2FAPCFS8jPFwCBHMRdGEWIKuBBt52I6P0HDx6OGju+gFJbEyxh3ngI4x0ODuaIT42DeB2IpeEIGaTXoiu6hHnewllI67WIgfwHQsBessMCR8JXCP6HonsBFFACLKAAYUCQjl3finCFKbZc3jiHxV0Iju3YgfiBc9ADzbXcQRCBOUAGZFkfe0utAz61dSMBUCiEQHDMCG7eMzhbiKrggCLMgcACTXokMqGGishJStVjihhijAhkKwkDSCXRf8DajaiF5rSXQv++YPjzJ7g94X8QCFdEhIuQ5MLh4Yn4V46wYMWbiGxYiCAOg4VQ20eCKBR4AQq4gUEA1n9YXPVdAXODXN5w0Dalh/yliDPVkAShhxowt0EYiEG4AUGgtFWIuwSGqS4bO2SoSTJA3dil4zNQ4hdQgkbF3YGkABd0Qex1xaRdq3LWjUYohn9I5SEG0lC+CNotnEOEiBNuZN4Y5YHI4YXo5NFarrD9h0euCBXeDR/eO4gS6L+wrkiiV4t4JKUE6H/QgX94gRcghBvAAVfIhATRgzWFhRXo6GNOgi+uYoqABXoQhiv+2JTmiP0l5jXtqX8IGALYOFBQLLhDu4qdSDu1wG7/+orT3c/9xObtdcxBJmhEheR/6GSO0Ne/eOiBEwjmaGSBeGqEqOcmAwSshAgYBliLuOSFSGWLGOWX/oeXTuWvBpEwqIOBMOuBUNumFgt3FotUsIiIhgjeo+sfhmUcMDeNzdiM/WJXMN9/qIBz4NUK+GJiRoiSXodm0GLSQghfCQ4s3pD+dYUVEIRdJIRnwABxcAK/jE1kuAI8nVY8JW0szIMrAMMwNJWqxmSISGcpJlvdyGeEEGuCZu2/EAe4FiSkTOvhuF0rKTasHojqVDoe9oXb/gdBQIi7hm2MeO2Do4i0Vm5cXAgWxggZbAS4dWuIQISxxU59hmVXaFO6lAI9/1gBV+jfhahlWgZWw14HlKbEf2hshADmicDii5CCFTDmLUhUhEjlf70BJ7gCERCBPJgDRvBsQi1LBfdsslTwDt013X1kcoCI3kaI10ZusSiI6aaIRx7qjqDkfyiGXxiI574aE+eNh9akDKcI7MMIfxYLo/RnGK/OirjOpf6HTf6q6voHa9g7Gbxq4WaOMKCAKV4BPRAGYViBcJDlU5FviIjvgYjv+abLCKLETCDmE6AJ/07ril4IfnaF0YpdFBCC7iUHcqgDcjgDcgiEMwiEp27ogXBx5RaEMFBugXjtYigGFoeI7LSuT0aI+QP0gZi97R6IqeYI6/ZRfdJMcfjtl/8W64WY6t9mDjiocU/tCB+niEsw9OUSchjniIfGVBzXDVCvCKRUBYjY7jDAgHCwAfntB2pYAUps7Cq3iAShxPo+347Vdfr+hyQYhHXIhBUQAoCmcP+uXdr+ByPcAhpAhEeuBWgH6Ovs0SM+6rkeiGwoBu/mjbHVdD8UbkT/54VAcUe+cElHCHfo7cu+iEh/w3JvntuldIxY64Xg8OVIOt7Q8X9AB31K9X8Q8uu7d2vQc4auCN2eYRBxBzIQAWpwAlfoBgjEdSdfbyn3dcdeXI69b4zgVSlv7HH8EEqc9bvIBG+ACA43wlyGCFowZWt4ZFpw+VpwxaKL6F3ECB2oBW3/RwgSD45KbYR/t4hi8PFi6HSL4PaJcPEKT/aNKGFa2PZ/LvrgQMqj7whbD6BLj+E1WAMrmWrs4/mqp4hGyIaAtwigZ+6BSHV4D440kAZ7cXpaAGglIANhoYZwEFmI2Hjd4Fhbp0tnuO+8/wsnTtN1CIFQTlyEEATdRvjXroXX3mQaIHVMFoLETdynlspGoHqxaARrwGpNR4ikp+uFnoh5txKV5/rr5HagN6JM+IfDHw6jhH2EaAAZpghuGAgdP4FNVn2EkOsAAoSxry6yRwist/qBgPl/yIZ/3/eBOPuNiNc0iP2OuAa0N+V/oAV0cAf4JQMzKFaEuItfdnKL+H6L/x8IutRNx0ZfjEAVW3biChh2Z+cNVWh5hDD5WvBupNRXuhZ3RMgGgKAF6F+jf0r+IUyocCHCWv8ADVSoiqFCaxQv/luhEFJCdBgNfvxHQeGWkP9oJRQihCINjBb/0WiZ8JfJkglPmMxpEk5CngjX/AP6cSLCCDlXIkSi0ySgbBAf5tTF0aS1bB8zLc2KkVucf6myocNwxQnCEFgVCrt47uO6hBUquNWatW23hGmRIMKp8ODFMAiJNkJ5ciGif4UdNvyH9J+OmwT/eUS4GKFNuR/1WsYYkfHSyksjN2ZYi9bLVBcL/zvhi1bBixgSTs0st0HmiKgnskKY+99uk6gXnv8NiQ4QujibP/bOCQjRxImIEMmkKEg2Q9MT07CKAy5OCCdkzYSr+xGuybaWyf9Dv7RCkkFpEbbNlHeB3skJPSO8tvClQpoSiSr1jxSNNYYSa//op5V/UGUV0XGufWQVIET9E6Bl0V2kym8YpZJgQoBM5RBNiOUEiV4mUjdbigklt9R7CL0YElFdrUiRf6oYpZAmDG2SX4rSYIdQV3Bs4t0/NiAknl01/mNeQhYypJ5WwqygkVsr4LBFbAhJoVxC1qgykFU4IkLTL4JRCBOTCC2oFWYreqTfg9SludCDOixgUhwTbfkPTYJ9ZKFpkPyQmVBrMuSTV6qYhpA0/zyaUJf/Mipk30eRmXSoZVPVqZOiWrGSxj9w8EAGO38kZIMZmdQV3EJ6xIjoQrFKSVEFNayQRELx/WMGEs3kmJqlF7Xm1D/NbYQQphRJseGxcnWKUbBC/sNNjap4mNlk0WpF4z9dDYQSURFwSxEPHPHA0LTO6JYQULTJmlOj7VKaLEK1IvQmOAilEtG+WqXLJr+QLTTvKVwuJSpGmgr1aDRwRNPNqQn98Yeq/9SQhKsI6brkRbF+9CLI/4yckB7mwVVBlf/ooVASK1CzApQ66XdNcZF1lQpR85o270dyLjTsX2yqUu7PCA40kLdCK9ShzxROS5F9eS60rEQ5eetjQlGnGEEz/33u5hO88MaLkS4K28GbnswqhG9CcfT7razZMkR1wp/qtAa7iixkyz/U2JBExiGt46RC5hm+osgXVdBWx/A5rpErFHCtE6boROYztVkPnEpXeyI0Z4ZyHayQwghZ69G/ZTM02aRrnh6S5pkVCttHtJHNOkJn/5NGNAjBEWmjERzc50LNXFQ6Qj/osrpsPMUukS5ysavsQnBo+tEa34QDBkbdDJ6QkromkYQZyTAC3+Mfkyzb4iH/o6sw5tEDS0auZALJ7FsptF1CpuWGFanIjbUuErCEFDAr6DIN5yjCkVMcMF4TqdyT0IMeZ1BQLtyY3j9+V7CypStd/kgFLoKnO/+dRCNIJUTIw06RighSpDfIA9Y/YpMK5Z0iOcXpnUlyB4c0nC4N++JgSGjIEFZML2uawh1D3hWDf/CNIWSpwcYWoqtuRDEh7LDFAnpkkh5tYh01UJJlRqYrL/4Di4ywgStWAAtXCAMXH3EGuxgYkunhcWAKqd3+PoK8GIIjN7xTWIu8wsOQVE9Sa7LbP5DnjNc1Kg7Wmt6+/kVEezXKg7r4lPIw0gwpsOuPHrwILuT4DzmW8oRaGWXaOpiQU7hwIdODgymXNy1IHKx0uYnU20KlkOwhZGw9iQYv48BBGtUSF8ozXrvyGBSFMJEhDSiS3xQSDiesoIoX0ZUT8kGKhfT/wgbVRCPHEtKxdXTDFeEQRslC8rj1XaQX7MDfP1yBvFP8oE/TEqTaugIOUU1PGqz4nSb5VajYpCuSfmxkDfnJm93kZn9y7CRGePmPDMpFc14z27eMacx/6CJr+ksID6I2yjvmSzZyfARLVSkXnkwDXq1kIS5+J9BTZqWWp/yUIE+alYctJHZ28ClyKALM3AWlASHI4j9sEYJ/hCdx4sPICs7Xi14gBKtZVQgZEdKyf9ADZlbSyfrWkQQntcWsVurFN5ORDGrUgB5t/EEq/IFDQ+pGF5dMCNr+MVM7RA+ACDlFEonYR4RwBDvRMCXeMALY6QH1IodFlNds2MFCnq4rHKI6WABzyFeE2AEOPNnNYnMjR6L+4wc5Uq0/AgIAIfkEBQoA/wAsAAAAAPQBGQFACP8A/wkcSLCgQYINDiosCGfhv28DGx2sV7BemoFfHBK8pLGjx48El4EcKVDZCIUvSKpc6TChPZYwWbJY8nFAzJsElRw8c1DAwDX/gOJU+eMfgpUTGBTk8M8FSGsCUw1VCDThzWNTFd7LSlBGQaBgV3ICCTbOLpaYNIYSiIokxK0LgXrjSrdjiTJ18448+U9LkZvRbgr9iEJgDyZ79sBUMXXaGkADl036N3mo1KwS9Eb+B8SrZrIw8XAlMvBFHHT/FhgMtGNHNUyTYleb9Lq1BQtRBnLhEkrBwSIsPgt36OBf8eHIkytkaupf83+ycCoFWW5ZOYODh/oUmF35Shmevf//TD7hn4rrA72IP6hs4JQZT/7lQh4+o8Ly09fHLFLr4BWQ9gmU2UAeeNfcc118FF5e18AB1DQDsSIQAANR+FEcBHVHVyQCbRfUPxAOFMBC8f1TgH4CPeLQIQ55SBAbT6gg0kqYACCAT5Moc8x16P3TI0vteeRFNQBU4wYbGzT1T4EoNunkPxKUt9J0Tq1Hw1wKVZkcRQZtB5lwXy70kkANKefbPwlM1YFCogGAyQitsPAAkFj9E6RAk/m0HYWYYFUnSX/+OZAy6hX040AWsLgITjAA8aRGTP1DmkYXXPAoUC9ld+CjBJ2pEDdvLERLmQOR6lEaHBYE0VBSepSqQGOC/7Smd3At5MdAckz6kir/ABBILDsM+s+cAhGb3gh8/GPJP8EKNGNB1okUbUnPjvRAe8oYa6dD1ymjzDJ3/rMdIVwIZNVCPHA6lYoLMRFcTCcsZI5GYWUXqUcnFrRBklO1pdE9tAyUw0Gm3uQTIKtmtcVAXJKESaHqjtTCmnA0oIsvPTA77EcjdGLAP4HAhEk14RbLbUHIBjMFQUGWbNB1xlL4Bjm/aKhQGUwI5JkF/7wB1UFKPXdrxCQNI1A7GulkEL/0fkgX0x0lQtAdBc1RkDqaFbBgiyBqxq5BI371T0Nhc7pVrTT8U4JBQ9v0DyT/oGDMyh/NqcY/yZZk0BQwu//so3sjBDPfeQUFMoNA5ZQTuCEDUdHJCNepwcfdAnXyjwEGoBHMy5yHqovNBW1NtHAiaDD66R45+k/AqKvkIugu/jOrQK2uF9wFlBxO0AhqBMKYCny5p5K2GVexA7JUCIRGFWj8gwYVVAwBTBVVBK9Q8skTFD0wyh80hECFcE/QDLmMwPfGiI/AWiAh9yzQGGV+TdC7yEEU4keLOoSLJx4x+Y8PC7nfP2o3EtCtpBLDSdNNXnIuh4QlG73yCAgG8oG6AOBnHvmLTAQChLLdZG0FKc8+yvcPK1BOBZSbAQj/MYURlMB6dJuBJarQPu714RaKAAb3FCEJSdzihwO5xT//miC97D1PIFWgQhX+MYQhNEGIIRBIE/4hvn9ETyO3kAT0LpeBIAShFSgTSPYGssSGQCQhcOCIfgTRupWYQCBWayNOIhCToQmkggpxhHUW0pCU/AMGAykAiwryRoF04Th1SQvqpDSLWfyDFzOYAV+CEQwqWGIb/4jBM2LxjxE8zxBU4B0LB5IscMSgD6MIB0jsYYcFdCMEo0DlJhawgBjE4B92EIgdeKCLzw0ECh7Bxj8YAYYhCvFjAtncDoJhuSAMJBiaQ8MMDGEJKqAgDUKZRn8EogWQLKI5bFhIKIxWF6bcayoA1I/UNMIzgijGIOTUiB2Hgpd/TDArKgjSoQy4/5BCni5vC3nFP+AxEEQ6hH85+4ellDIdBuyGEIQYAV9m4EwmkuAftvhHFrQXhGCY73dDdIgdJEQQVuBiPTwQhCQKYomKZuByY7Qi9GbAt3LsIAoQ3KZBaqSR54xFIQegizn/US4B4iSdjyLpQd6pl1IYx6moW4M0JAISBxg0JhDsCdEsNRAGnFMgZyBHLEbAGIIg8yAGOMI/CjGQdMWABu5whxD+odSb4KKuLGEFK3hAAXEAIwgZyMD3KlpRg3zMAFQIAvQ8+oByKKMENHnS1+QnR83ooiB/qadCovMRN3REFDhZw8JiEtmBWAUqVFuIFbhqHIW4gyDlMkpHLCSQWv8IIEAjKZFGoHqQsKwqoR3RBTlykYOT6PByyD2rupR6UpAgQ4wxOawXE9sKyJVjEi3c1j/CVNnuqkuD3h3IRRzzj4topKzC0dZAmpUV0OLkOQQhRCpo0INcANSKVViWIUB5EO6dtbDH/QgPcqmLAf+jwJdtXRAMsODpUqG6iZvEDl7gi4opBL4DOcFZ9MKvDWDYIblRCT9hMmKVjACPP+WUVSBBgPywpAe8KhVqWOLeJzUAgx4J6j94SyKBsNYjnIyFIQzAuIGkgIkDGQIGivKOgQhTIHooyArMkBdxNOmwmDOAJRAbhP3yIRCTAMAkAoECcChhABNoFYbhoAPkbCD/xQvhKgJXUiuiDSwmuC1IAgj6jxor5McaGUs4BXIUjySUdQoSDhOAOxDwfoSqAqEfUHGSv4XsIMgCGUGRzToECjTDH1FWSKjPsZApfka5ODmyQFQ9EMylAHNe9KLmdiDmBzyhBS04CCLGlhwthVddaaHtcM5ZaYNs+B8JnXNMrJCcv8xHZ1wBINJgYornQG0gIXsBCpRQBT7wZQj/kaJKmpuXdBWkD8VkhEeOzOqPfK8gBhiCAV79agYzWGXlqIYKKsGFXHtkDiJQ1301EquhNMsXTvt1R17gx54q/CZP8GxHKjMUOv5Ds3SxeCYJYm6D+EMguAi1XirQkY9rJgVD/0iBylP+anlbQpJTUEMr9iGQoRHCvP8QjUeUDZIk7esfchiOpIm2ttI+fCSi812+PvOGYLXTIy4eiBqHA4MnLBpnZeAkQT48EE6slC7kboZAiqLx7n7vpe/+x0sJkoEUtP3tble5IUpghRLwYh+7GaAfPDGNejQgFQJopyhM9w/CH50k084LEKxXVYKo7iYY10j+NjBojej2HzxnL3qFOpTmRF0g1xDIqz5ieI3k4gkXuDoLDuFVXsTCDxzgBBfcgBsVRCEQxgj3Sm5JEt5rxBmpAX5q3teNf/RhIIrwzhA2KpAsBDYDzn9+YDsRjJlzgA2zYEBSBiCIiq0hDbtwg//6cvAEaMQzK8X2SHk0oOO6BDXxbUzJgFjC7OQwGiYKPIi/62IKBkznRgFQDByCJRDTTytRKUwAAx3gUNrACwLRCjMAgXwQCy3AC63AB60gDnkQApuAHOxgEKrUDX0QArYABr3wCQLxB//QDck3EGAwBsBXfFPxUhtFgwuxDVkgD1mAgzqYBc7XCbnAC5aQN2WgQiMgSSNgBbwjUepjDNswD8OADwORDlPxdCBzeC9CQHjwBcL2KJXRTR1hCpQnEGzgNlZYEJVQAAjEc0NxVQtxhlf4EZUHZwAYAAEAAF7wAA9ACZQwAgHgDS+AAKigAJ7yD/5EEh3AAf7HBQzABqv/IA/bsA9BEIGtUIlHxlYaoRosQVkF4Q9NJhDr4AQCAQZgoIn+oCJf8wl/4AxPBhOYWBCvKBDy8A9qNYtqdYtZcATycARHsA98yAsWaAiViIHUZAD7EFhxNwTykA7F4WcGAQJvYAE7II3SSDcCMXkFYY0sUYjCYYWmUHn/UGnstRBrE3lckR8YEkFdOBACsI7ph4UqAY4FYSM3sgNAMAUPMAKUUAZWgIRqcIS8MAur0BsK4AKeYCMAkJAAsAMqgHq5cAEPWQlPwAIqwAIS0AMqAIzCeIHBIENqt1YfIQX/IJIGIXxeMxAn9Yn/oJImlxfMxw8DAZMwKRBt8A9tIAbI/3AE2wA9LyUG/yAGbXAEYnAEQXkEWdAGoBAPXSAKDsCU49CUDhAKBVAp5WMBb8AaUxALXMALfiBpLrApMAF/IMEJTAFnB1F6BPF0cDg678gVS6cQWvcPl+cQY9GWHSEH62QQFNKFP2YpIUYI//B5AhEqB5EDU5AD12IIfpV2rQYMmjMDHYkGrdAJnSCEQliBlmkJmckLlGAJlJALVCAPkFgQzKccJLcSKukQJhkTvEiLCuGTz0UQsdkGNUmTyJAFBpALmumLwLgPs8AM+8AMXLANXLAPvNACfAiErZALhpALueB2R8APq9BJIxALucAFzKAN/yCPGqMXkvZVyGGFDf8nEHPJFYX2ETi3Evc0NQUBSDhxHOMwOpIWIAXCD2tHEEe2dmx1kwUxnRoBATYJi/DoEWTwD6o0FbV5EAmqERdVEDW5oALhkxL6k2olBhDQBhDAD/yAcimQC/M0Fe41KR6BAIL5EevZnQthH+M5oCPBAhLHogdBmCPhAgUyFqGQB0a5fNBHi7PokwYBoB0Rm1yBBCRRdo8yBgbqEUAqEEs6FavQpP+ADA8qpciQochgPDLqEHkmHOfZEcESKic6EvfUPjBqEDpnEDBANUNnKwYRYv9wCDiAEx4UaQcRdDGxYWYpWwIBCIAQeoDQCJGAB+SyCsiADNIJAU9KAoq6EED/OpsDoVax6JoEAUwfgaQgYXE24BC3tJp0oW4BiiIkAAGhCgGkigx0wAUhUzYIBxNnAQMv6hBvcBZ4EKvrMQBuEzEUsBJrEBj/sE0gECB10BETxD/PEAU94KY4sRYCoawHgQX/AGkLEWJnMXUDcQPIARlZVRAbJqi5KhAEIAcE8A9noARngAFVIAniMJyrcAVPSqhrxVZm4ArhsAU1kATCUAFESnJOYKlEmhewMBKDIBDh0A+Y5BHIAJQJWpOkOhAX1aAE0bAEAQr/ILESy7CgQAJ5AAoZ2wsaSwK9gLF0IAp5EHDmURoDMYAHIaJI9A+XcGwsu6pNQgjoJRp44As0/ysQEzRBKyocGIBHKvElYUIqDXQQojF12dAIxYAS/7CiCPcLI4GsMBFjCpG0IzF1K1oYchoR1oAlAoEBgAmY/6AENyACoRAKqzCyhLquV4ADriAM/3AOpykQzZAEC4E1A/GvMKEHzRC3B0EPK/APAasQV0CUBuGTNVmlVcqkoHAFt7ALgVAFhXC2q0ACkyuqkzu5JHCxoLC5GMu5edC5dBC6/DAENCQQorgkBoEDzgoSqysQ3dokOHC6obESl4C1MRGsbPQPmvAZ6agQGMJdAmG7BdEfRnoQYfAPMJsVOBYxCfYPqcKnwLu0GpG8A6E0rnADrpAJ/6AHFUByK+AKK/8QZXxLcnogckmQBN2rEJw6EKR2EM3gDHsrEM5wDu37D/haAwKhBMawCoRKlEBpoRiKoaSKof8AoA0aqmPgC76wCwq8C2egA2cAAmeAAkiKtTqBBRiAwVjQugVBvQuhE21WW5HwKhwyVwMRrGGwulTrEHEqEC0cUh+MARrxwgRRoAThC2Wzws1KF1QmED0sECY8EKMlEH87EIJAkiBxDw2wBt9XJrlUEA0wDXAQDekJQWmjEEaqNLqru1psxAvxWgcRY5ABGTOWiQ5RC7/QH4gWE737EXBDA22mAzqACKEnELRArf8wCmYgAv1gBpmQBOvwEYEMigexDqRGcnFbv/X/qxAimcgFUQOusA56kASuIATUmrsDEQ5m4AQiIAJ58Ml58AodmweiegWh+snxoAC5GsL/kDZXzEaCQA5g9Q+79g9O6xAHqhFSOxBB3BHZ+g8yHLj/YK0Dsca9qhCyXAeYPMzVOhCvOxKYLMsDscurEy+sHLyXgMeuMBDbTBAnQEfxQqRuaxCaSGI3sWuqULwF0a9IXBDlTBI/Q80rcct2rBGjJQhbgMm7W8cfERjNaxCXlQpwsABO8IFEPBD4SxD0MBIkN8j/sA4d2IEd4dAEwbeFDMl0O8h0Sw3ZK5I6YMLusAX0qhCQoQq0YNKqwCsBQ8+0TBC1/A9z1a//0GbG//wPoyXDNl0Q8fIPdKTO/8DPDgEVgFDTCrEAcDPN/2DStgzEwwfTByHDRRzGP4NoJ83U/9Cv/corKY3UBXHFq7NdQ1EUIzkQ0hANvJoXYREUDYEL6UnWAwE3Yj0QxRsBzlABJEmkMq0QMRYHl+ERu/oP0iAVR91xbXzUUeEQ7awQDdAwBBEYDREiDbAJTtCCA5GpTrACK5DQBFF8dPsPSdANm9DZcStynq0QFD0VSYDZ4ywQ9voPwvC3mE0NeW2/A2HR4CDPA3FLcHNLvCfYb60SvUwQkKDb4KARkBABHScQaXBZCQYIfb0Sz10QiODTA4EEhg0TvgfYB7bdAoHbT/+S1kNRKw1hKoGRS81FbieFC9GQMB8X1y3Zkm4tDf/ADSRlVLwmNqWCSw0RB7rADTihC9KAVw70Dw0wBmaQUQJhC4oQDpr9ETJYEPkgEL1ACgNBCqTQC8nwwwaRBPQwCOC72jjRDaKYDP+QD+xgBtTwD3/bDd+bCXsFCT9QFP4QAT8QAcftEObVXHbwz/9gbuQmEMw9FXiVS7kUGLiwBo5x1gORjjxw3cE1EKmQCsl9Ur59EEVRFI/Aq7gg3wIR4ApxCsmdYHbAq1/z4wMB4KfwD2In1woR3cJRMB+BFYAA3uXVZpnxeBshIs6b32kJEkNbEEaHIucyfwIRAIDg30r//hFrwY3I8SAfUS3JMXSbJ0d2ahA8cRCjV6YFpRxtzRW/DMV0cS5nahD2PRDEsnmicxMe4GtU8SEJU7UOoQBWw+h+nXBEKxBcmyH/sBWJ3i8CQesksUJ14VQ8BhMlel5zShKl/g/8cogLgQtLpBHZ7RDhhAqc1X4swVCBqdfC0hHL/qwaMSJwzinXgeeaPhKJkJeVwAcscD50UYAHMY4CIeze4WgGEVt0UWJDocNWPRISYO7Lqhzh1Bz+8j//IJaK9y8oOeDcUegHkRB/PhCprhCB8UAjkewGMfFk8g/2PhTZAYYjsY4DMQerwAm0tyMTNxAUpxKBshJD8g/VYB5P/7BOSpGn5y5HWkDoHpEQX8OdwyFxXk0XZdIwqpARFiLyH6HvDpFaBDHu+O3wDnEiGo9/wG4QhJ6XKnvYRysuEk8J2hgTsAEbLDMQh1IQ8M4eKlEZPcAFb6YkMDH1nMIUx04QgDYcX6nYyYFUesHlCjEqBfHtCpHpT88VuF3cmLIes63wIFEAKZEQqlA2PRALPdJYaL8xczIDLEAy12IoLe8jhVIOdQL6HqGQCDkQu3Aj/5C0qv8PdmiHxRA2IxIAjQCzBCDgN28QBZcX3n2NAw7ekWKXHrEBBf8Rs4LxOOH0Vn8QbYz6DV8XSj8Ss9PoCbf7BxENvGIMPTAFK1P2LP9zHSOQPYxHENw/FN1CENpyHSvjN6Z+HTE/EHcQrh8xcBiRHC/BiZrB2CCR2ARR8MMPEP8EDiRY0KDBAgZd/NvwD9pBiBElElwz0eLFg/YmJqo08Mm/HBhFDrQz0uRJlP8G+CEUrQErcj2mCASCMZbAmSkfYMJU7sHMclMsPCg3sKjAo/+CBkODxlCwoASVETRksVxRAP9A0KqIkcnBN9lSjr1oiuzAZgPbXawztmI9gScOnS3Y0KQbPHQFShhIS68Ago3g/Gvwr6teuBJLHgSEcYJei9/+SRZIY2CuRIly5cKCJQwWgb90KemxI+c/NTgPPhDI57TFKcH+jSg6ZUT/MENoqogTt6NgINn/dv0zRkX3PyoDgY0Y8e9pxCqzc05NyppotR09xgw2HLHEv4+QL3YRf3FPRB/l1a9nr7dixVTtTwqwdthgpIIlEqa08M8v5DIG4sKPXFL7RwWDUhuBjwMNmunBgZoTiLWBqrhFtuQyRIOKDK4YYiBJqHgtImA+/AeMQhQpJDk0DJKkoBeTCyYYS3KxJBY1TnuQhX+myElCX7pqoCQE5TNIFCOTZC8RJdmD4R8e6eqqq6QgGuyFs+xDKQCDlhiIySbLI4AcHBX8JxcJCVIjlibIyqMXDyUhQxJJmmjillsiKoSMK0Rip4lw6PzQxH9aRO0f2YBJ/8EANAyw5B8AAkFBF8IgCkmg5r74hxuIOEEpvfRS4iDMgbRchCDy4OnCBIm0JNWgFl496DGBOI0IiGUIKqwi7lIi759pZJVIhol+1YsBlXaz0RIDeDFgoD6qmPFRKqpNc6BnJApnoEIOsoOVf1j5Fpd/cOHBDh4oXUwgHkRyxYwVxtjknxhikEScCIMJAjmCqAgihQxwKqeaap6xbLJiUDrVLIju+GeYA8QbVaBRGfBEWIwxCbMUjA+qKaJoOv4HnX8AMygvsg6m66uvDHpsAi48CaOHawkCxiJxbpotluj6OEkXcAuitDxdFmjCxCCCuDkFfgsygIqb/wmCimBoq/9GGRYsmMkKgRwRSFOJ7Joo4pM0MghZZNtbaywNiBb5bYJqLqgx+bj4ID6BgsWoCPY4dkC9EwiJ5dKC9oV7IHITR/wgcg3SJYZ/jng2apH2DeLpqammrRwvRpghh5o+bqyww0uHDJKBOviHiFf5OqiUcf5Bsm2U0ihVoFNPahkEsh4aaeL5/tG4PI4H+tugiiSbBhGX/8mdoDD+QSEXPpqzhPJnbf7nZspNf/Vy8IPYEA2rJ5lCgjcwYoOkf/rz/v2ztKArK/hFqkhvg4h9G2X22kbSpD10JCIR+McLevCPGQRHIIZgmosoEI42CYQCAxHHi1ACLgz+Y2hC06DI9mX/AANcDhghtES1WmE1ALwBBOC6R0Fyx7B/hAxLFtGGSdZHEBhGRIACycVFCOg9/GQjEvwjHOEwcgmBeAMix/sH7VCCB/y4EHhjoQxE9uM+Iy1BbiH52ECsgbx/gG0gvIMI2f6HkrTdkCB5iYJAKNGKGchtCCAUxxYe8YhTVOAgejiLLUyyAhxITVYgJCTmnBKIckwCANVggRt44YeBMCCH9ZPPHIq3HiUOxGSQycoxCkIBBJDlgGOJA0TO84/v/KMWlBSIxsKDyolQJlfqSeU/WobDifSAFwPhw6MGYqJMCGMgNSCIGc7SpgiOJJBkaaBImPZMAyyqkMDwVyumMIly/yjjJgR4m9huV8WDnId1rGySxjxJzlbkJyVcg4yrLKK/kdAPImsbyS0hcrGBIAgFCyCDE/6xAIH88CTv+Mcj/LEJKQgEcuTESAOH4NAULEqiILSEJUYwhaA8YRYRYR5B6EmXh6ACY75jKPyaM0WMvPJwmLBA+p4okDg8YiKTEM8TysCEMpShlpL8xyQbhJEf/uAi/sBF44R5ioDSJaE/JGjHPpSBFDz0oRF9qAGqpoYRUGIfsYKkQKJRjzWkQgAzVA9J/+Gpi1RCgAwYhkkOsVGBoPUiPeSkReT5PkiidK7/2OFAfENOWv1DrwW5hkR+EZEzRuQCTMApTmFABAZwAf+uPR1IIP4RhSpcAQMmIeBCU+JZ9XRDPgETSMAycFqonjYLAIPqU7I6i238gwETmMAA6gAHsOoiALxLhxwQIIsDOJEuqBMJJQaSjlCV9CIBSkmRIJI2iHSRWPBkT18JEgjnQle5EfGCRIwlkguEVwYlSAQXuMCLWDBoBv/gQytawAv4fmgVZEgJQFPyiYLgF78HMYJA+isQUhjhvwMZ8FkykIWBIJggCj5wg7PQ4AwYwhC80AYHKswMLuzDD7xwQyymkKMRqEEFamABF2QhCnwM5LsF8Usq3KkXsrUtdgs5ScQ+Wh6N5eWu4iHrRJRwkFmKRK4C+etF0lmeBKyYPRz/kGt/BBCAAEQCygDwQpX/4QWa0o0uT1gseTnAgFloYxX7eJQxZhAEXhiiFWuWcAryoB5sSCTOjLOFgAXyB2dI5h7OsME//msEMIBhDOvpljz+UQgFCyS2/8iCPLKAaEdv48GdoEQLqNDe9s4AjnEsgedmYAlepAAYXJjDMGYnu8vs5zcowaJIEhs2u3gzTHgQo6x0MJAdG6TWAmHYIswCQzISpNUeEdY4B/IGl0JklAUZsvAEIgBoA2AZV+PDegOxmW24YBWhUIACEuDtBITiDgAQAABSyFKBXECA6n4CCxLxZQbEmwucmAUl+FBtOFJhCIUeiTP+IVD1ENQf73jH/yOwYdB/zJkgCidIu8wgWiWJQSBHEMMRjpACKljC0PywuKHl4WhIZ6AQ+34zQS5ZgPA+QQItDYRpdtDyQIzADbx2QbOLbJALiGd9nlIjQZI7kWFLxLIC6TFZAsC/s01kkwbJJGRi0cMe5twiDOPAIrSbEgJgMSvVEMlgk/3sf2hhCkCYQg4oMQM0VBQNVQvxDKzAHBbMIBeU4EUi7J2LWCSCFy2ge6X3PgsM84LSlG5FLmgk8oAlmqGNs8i8DmLflBwhcv9owxH4MZA2SFwgyBiIGNrAj21Q0xL84AcySi8GZBwBGVfgggIc0AVRdOH145C9CVzwhHtTwu/AqEos9v/Bi0BojAsC6bnIntexr1D3VXdtRGAuQgiL5FzVFvHUYE0uECb+o6sGWfpAaknsi9xcIG2UirkPgYwMbIO0hDJCVAdi6H9w/h+rQAYEkEH/1JO+DfPn/P7FoPn18Lf1YDi6gDyMkLz9O4gEhIB/YMAGjIj9awNkkIdtSAFxsARx0L1O6AQJM4SKApiP+wd5QAYxgAAIYIYSygVeoIREsIRtYAZOuLqUuKSTYIBm2y6RCCWCWCa6kIOIGA7ICKyIyL4wGQCB4KaJMCKCCIVVAAVEIy3SKgj5EwgHHIgqfBUDxMGTcEAHJIGB8ELx2D/OkzzK87z6Q4Y2OC1xGLp/0MH/jjFCk2ip9Am2McIINvSeTYoiO+AO27mI4fiCr8ufk4DDZTsIeBCIUJAILhnEgcCB7ROJL4C+gXDDgbiESCgGCti3fRM5BGRAMATDfwBF8XgzdxCJfhAJAUyJVNSLCDSILgwTE2wDCJDF+1sFLkgfwEC6iUAZlwq28FAAk6BDutBFjCAjYRQIldLCg8gLYtSZsXAYuogiiUABahQIH7RGfLlGO5SIGzCIxlCFgrAAEACBXQgEAmhCOgAFOiABEoCAdnzHWJzFyqu8I8iCI5CHeiRDiNisiRAC+aAGicgEgRgFjNAEixBFkQCFgVDIgyABUHBIdiQBRmBHCEgHTiCE/6ADOyC0xosgRlaSRG1UxpS4tYlAAbqgAEm8CDj8B276ANBwvoLYhV4sHZLpPiQSCE/Agg/4AALgSZ48AxSgAaGkgUvwBRTAAgpIgnP4h6UciKZ0yn+gB2JagX8QgYFAgpMYBJGABVj4h660CGroE4EAQAhswFk0QRNsx7R0R3eMSLd8SLiEyLgEBbokgTwAhbu8y1eIh1dYhX8Qy4EoOoNYRIwYDl9gDx9kHWOzSqs0iJQciLzYpEsIA25CwjDhx+gZCPoqD2mgm0xqvoMAzYE4zMAkix9rxH/gwdQUCH5Uj8dMkj40iC8SCH8UCHIgCJIkTeHYhTOwLJPcrBughv8a0AM9aoYkIAiurAFXcIV/0Mp/YM6JoAd6qAA98rdVbIZVHAhnwE6BSIvurIB1oEqBMAcRsDjTSz0JlMD4K4gEjD9QWIVn8IVdkE/5LMp/OAMsiQJy0M8zAEolqAMKCFDo+wCUBI1aWERf0E2I8EEdICsQeLKLwABCmCBVkpW2GAgPmESCeIEH/QfCvIgPuM9tLJ0qWgPSkYiQkc2IUJm38Qtr0DKTWCVVktE/sghAgNGIUAKSvIjb/AcKCE5qMANh0COmHIunLAgiNYjslIi0qACqFIYVCIFaIE1yIIBCyINVoD/7Q0u2hMd3rL/3dIcEHbRB+zEdQAHSNMnMLAj/+6yFYqDRk1ilxpjNgrhQFqtQg2hNg+jRf9BNGbWstljTgbDMf+jGbowIOH3TfzhNgrBTkfgxJSBKgjjUgXCFZCKIhNqCf9BUgeBUlGghgeAOLXkPglgX//gFRDgBGjiBfzisiPBHf8RKgmDVE6hNiLBVgrAGWrAGVbgGcLwIW4mIxvALQKAFFm2Swuqof/uHUhqIX4iDNvGnhxPI9ViHgbBWgcDWsUjSFRiE4xSIFXAFWzXITsUA8TSILdABRECEKZ3SPnVXy7g1HbAMy4BTRlUCf/wPWtjXjjpXjCDWXI0IVu2LhImICaLQf2DVjvoPiBCEgbi1ELAIZZ0IgyTX/4tgWHkNjYtAqnZpF4FYRVn9h4RqJ5OIzV+FiAgYWZEtCMj5BVVgVT6yWFtVWYFABLw5CVZIBUjw2Ii42YGABJ89iZDBn4kIGVaAA4BShGKyAX8dCIgTJm0lCz4yCD6K2pHoVmHA1iQQJglyBfHc0X+o2LAdW38Ex5MVCJIBR78AR0hw1ZE4W4twW7eViIEtCLg1W7A1iPiA24MY2Cy8CHAsLIEQ3IKg2YEorJuND1tx2X9gnl9lWIIUSYkYjBQdiGkImn8QKqTyB6T6h/gAF579N++ECKRqVoJghTRghWio3F4RiDXgFYGwg9g0Xb0AB4FIA1NtlQaIATDoM4PwWv+Im4jgFYhe+Ad28COB4Np/SIJ1UN5/EKYk2NokCNdvNQnnLQjHo8p8IIVkEAGADNcVIK5llQhKuVmSEQjMjYgf6NyDSIWgFY9TOAVWOAVcOAU7oJSgKaVmFaqxEF+CiN+BsK+ESsX4BReg4RTTxRvQIgihohQ4IJdHgIOhAZf3/QdwEKiQLY8THYk1aF2IKAxpPFyKIAi+EQn+IVr7IYhjOCeCcJ2LWAYKkQ8ZkDq9SERZUSKZktyJeEQd7g5lfAxfGwi0koUlMjaCYNiz6D6T+FCDYOF/gIvDANsSLgguYeKCeLGB8OCB6C6JeJLbOYybxIgbhIjDSLbwkIEQHQv/kUoSOvXIw0mMMXLhsUhjJXmM4WtDifi+gYiE2NxgiZCGLKELGjYLNWoIIiabgfi5O1USP7bRiMDig9ikXBOIwngEOi0IaDyLYCFVgciLLpKIMQYjSBYJ+SkIYAzkRu7hgvBi5RJCi2BlgRi2VDYIh+WVED4IImQcPRWJUyK+giDijlFilIDjs8gKwNA6VU5hiQCTmYuIqTCIBCiINSYI1YkIDx6BHBgBCciaBB1HC3i5N6CBbACHOICDsNoW9VjjObCIWVaS46FBLSwMOGg6iGCVJkGrGyLiG2uPxjgGL1gGKxOPWx4IcMKITE5mZT4LJRSIaMYIMCkAN2iO9KGp/4OoBoq2aIPgnILwAmWYgh6AATCxCDpWkik+iJVE6LPIyJESFq7DiGnA0YOYhq4Q5lEuiC46aPa4FHhSPpS2iB6YCi5+m3JYEz6wp9VpEgkogkAsiAFw5e3aNbpwLlKZIhqTFScGIyrGCEBgYpg2CDeYrpOAi/O9iDXwhpIuiGSEiI0sD9gdiISYPolwY4JYBW0gAhaoEqQgCIqGjJZOiR2QO4E4BLhmKHvu6Xzai39waonIYSYrD1AxksK4hFwJMorQEpkanlZpDCueiMGWiDDuGDhQUIyY5kf+h17RY4vgH3b6h3VmAzd4Zow4J0y4aKMQllzxgilggbmQNdI27P/yWOqU6DGeylBUsGGBIKjDkClP8amxeAUfOABFJggZ6OzyKCxSLYwKFojsNpK8JWuC2Gz5OGWBEO+JkGOCKIBqPohLqDUO8IMowGuUAIBJwAQv4DqNFoigThLMtmgLOISec4EMHQmwdgzFVhIZfJ8AxwjrO4voZiiSgQu4CFasVg8sboQ10IjDgAMu+eT2wIE1juaGxojVpuZ/SGPsLhnA+IKQaLejiOGx4Dr6TgqMJggvgG/xgG1cax8/AJ5QPonPLogDT5I7HggjlggaZo+0qWpRdqFfIwuHhQxUoDHjNomaNggIbwAJFwi6qfKTaOfG4GSB2HBSWeckQZkveIL/i8omiaBsgVCG/D6ISaiGSeZiG4+IYziKY1AGFs6VO/+HZ77to4hzRcIEAkCA47sI/WGuf5hieoYbNxzy6BOIKGkP5v5iF6KY0ultlAAEDybmkQBvvejuieDy8sDVfwjxggDVf1B1iIgViTCGu7YO2H5mF/dz20AvZVDzgmBzZ6YQHIcI1lgGTBB24Zm2Y8CErFgkc3s2CB2IZk2DUlLNVZeIQuzhgj4IJugBlSaLSj8ILWnys2gI4RKZ1r0HD+YLvhFmWfF0ckL1EQbzkwABmqkOifARZwSyf+B1IymKX5cKglBzvAYBIriB7R4IvvVtyCiMdjYITZ+IHj8I19kA/7NoCFl7Gy0m34FogDWg3ZLpavVQd9Mh7yUn9YIAAQ9TCpH4NGAIhpyoc5THd5e/iKCYAYx6gH7387zGeeowCAvAAIATcFkxG1lBYYiAY1EniIZPkg0wK71w94KA0yahG3ZHeGEZjDQIhFhAJJHQJrpICo5GCn7H+YiY+aoIBt/4iTbPCT44eZEIBERY+I60hmsfiAVXLn/wJ7WQD1LNYbip9lcpAFiOiKWDd4jg6YkIAKiOiNwVCKMmY/Zg9YQ1bxLX7gZQBSxQgdfgcBzvaAmjDYjQkYKYiplgjSn4iSnYjNJP/YIoiqu4jabAlKPQkU8rITSYgRh2cWVYBmXY6/9a4HJFPwjIfxu54gCEvQgvFlwiFYW1aIfYgQhcCAPqtggtiX75YB0wwel/EHmUIBlSv/iCEE35kOrS9n4jcXqCYHXSeZISYIIjX1nXHQNjGBF/NwgVMITmYP1+j+GgGIFWAAg1D/4RDDTDkCEqBBcyJDji34iD/6osTMFnypRYDIP9Q0NwSMN/A0Mu3BEIHMmQMMqkbNmQgcuYMmfSlNmuJs6WbnLyJPni38+Uc/4NrWnh35SFtHrGjASHKdSQa2Q+YTghKlYa/1iUoNSKBZ9clFrw8sNroacRanjyaZl04ZRgrdCMCBQoGBoqaKoAA/mv3N+QwUYEC0aRIBVJQ6r/UOzUsfDCxAuBEVyL9J+jkOWqWajr618cXbpi/Iqx8CnW1P/qqV6Ii2GlhSx6sv72Tw7UqQR1y2jtu+cSCUsW1vr9D4/xnLp112zxz0/ynCxbjFBRU81bkgPX5oBLUIXGfxw9dlTYkW+hQv/+SLpM0DHilJKa3JJk4J95l+3N7wjWiYpaDSU1wgibAfCGQ/+k0kADoKX2AVMYLDRNTZwQxAFBrIT0Gkmz8cTaP5r8MwBTUzH3T29RsRGdcY/MZOI/17AIFYUENfgPILREkpwqv5XRGxfOJdJDdg2pkEMu3f1jXWUEaQEXHw8BBtE/t/wjiSTm5aUYlgT1EUIThYhT/5gh+DWkV2JZNNHQEFkGwaaVDUkiDhVVKGRACvf9o8w/T/4zw0MdSdXgPf/YgRxOMF3IlAYzOhpTAo9KShMIBA1XQkioEeQiTfWs0eMyMcEBSFCTpuRNAAKkJsFvgchEiYcxjcAHR+6JNEIuVbbH0BVgEGTLPyGE1AeXt9RZRV5UGDCEIvPdEmeVH/m1a0s8fMPDLcAAQ8UQGVD2ZqAElckQGsDw8gw4hbrEkgzD/VMpTb/EdMA/9Jr62w//rBgSPP90EdOJv21wL0FHuaTpQtDJ5GmPBE3iEiDw5lZTg7oB4g1DAezZ0CEE90TJZRj9QwZBgEJUpiEPWebQYe78Y/9DT2tGK2wIX/bxjzvd/LNADJuMsYC8M9kC7D9XkNyEJCksFEwgA1KhEBXAcGFJeMYQgsGCNeHBTUOLMEXvTT6kxgEnYUiqG24YLmRCTQHXBEBDexDUgccEA/FPqAzV+A+FEmNFxFVQaVw3TxNwoA0nGewjzj9v5kfQL008xEedes1ga0NpNITDQlekxAMPuvwjuuiGmt5aCCE8Syy1MwQywptvNoRGEAYYslkgOqzh4hoBFJETB2pb6DVJwxBkr2pqE04T27/BLVNRLnX86CWq3f2PF1PyzVTzBP27fEgpLvRZS93PxMRLDXFBCCHWYTfC0wxJYidDndT6T3exkPP/S9AELbAQK1jBoZDYAStjCEk4FlI60QyQXGZS2j9SkAF55IkKlqBCMKawmSlE4QRruEcxQuKulpiCICX0yR3+0SjjKA98LiTYKwhnMJHo7R+6icMLjcMSrbjEAb5ZHyEIVDJL/ENPBGGPESBogAwMARjGGEFSkgKtmmjoXqO5hV9IQhkzEUR2T0PDFKoxCZP8whpfYIifFqK5kHiNeCRJoQ/ENpMbyaSFyTFeDhcSgMFRiSCtkFQpfJjHkEijETkR5ExI5BI+MkRVeYwF+hiiqIVcxRNheCKTQrIrAxzhHyTwi3qARg4MGIMgz/hZTUT3GlzwABcCbKUA/9HAnrAC/xt2cIc4thiEDGRgIUGQXRERo6enYXAKO6jGDkYwm5UN8l43+cczoxLIGEoqV1g5YzNrkgZA/INVNUEkTlhTI7fpkSCYUMbvpOIaj9mRIEJwQw+UpC1fNu4fWySJzGKQigxFBxerrAmHWGEHXYzBPlnopT0XYkSXBIEKQeiEITToBWWMAFNOWgg3Xbi3bHKUILLoaEgYEDiCqKshLGGBkkLCDWswpRQz4YKCVrM9mqSzJcwRn0tc6lLjnCEVz4iFdWZgCcrcs4su5AFBVhnLlmioigv5A2KAiZP7GOCXvzQEGMsxCS+ooATYaYg9QnJCkJKVIUhtzSxykkaXiCIqzP8x20ImGZO2LARBTLkAKv5hvn+0tSUIyIkAMIa35Ihipy7RDQpqEoY06CAXJksoQe5D1MmA74A4KV1yqlpVKhiiFRLdDJFq4kbMlrW0LvnC9aByjCIUIZOMZIgoVhgVhOUkkuJjzRpoGxNo6JUkkPiHhEI6k2M0JJ15Mw44GRLWgF2AIRiCCQNG+49YdEKIBLGEAb6lrapCNjq6OKtpG6fZpyEEil6ohjJ6gKiW7OsfQvhHNCY1MJ4UIIfkTAkOw8uiqoSEQiBqSH3/EeB7eeEfz9sBi/pKE7oSZMD/sBBDEEGQnYTLMXdqyH2AWTujxocnotMQaTkaO80GARi/REP/yrQKgB2cARD3ffBCXtyQaOKEExuY73xjYs1/xEa/DXltSkZaEz4BmSHjYMoaf4MOG+ZQQymlSZIXUlKGuKolso1JJP8ht5n8hA8z6EQKPAKfyShNHAuwB4XU9Y5T/CMCSMiEK27AOWqlsplEvK5Ci0jihgbBEMHAjhcA8AUaaGoCE4DpP9zIkCiEhMYEeQL5arIB3rIBwjPpMU59nBziGvhRMq4Jo3fjEv4WTFLPW4gjQ2LXkBjyehaViYJbwuAt58QSf2zLWSpiAElQYBPf4NSkGGGDTBAkEyuAxSDCYYa66ckAzgaGAZTFWTQEYzOTqAYIdFAHOdDNuTVxNE8m/60vnGz51WTtQKla0p0n1ySjMfqHbn+TboIoWiZZnhBLYzJD45ygJpnEyT4b0qgrR2WsIenyQwjkGAhWhAJI+Ic/mgEVmbUGFjcgnLMzXtUgoKETgKoGALyQAwcjmiGfduGONf0owaYk1gwh9UK82RLi1dslzSUIpjSWhuKkJBGEG2GmkcsTWp/Q4FT+RxSsOZtW3JkgSiODOyTeED2QZKM5IZpLhLGQZf9moS7Bk8ah7dCnFcgLXIUnSfIlKRcQZGCKZHJIbr6QoCcnjik5ualOLUmo/Dsmll5INgiy5JZgk6NZ3jfdTWXuC3HAFDlmyAsMFggQECIXDxEqwwmyjf8cakLtm8gj2DW+8RSXwwss4IVzFvL2SeV1A3//dI97sgKcEHwhWskv+EKFiXthiA1eY0N7ZUJr1URqRqltMAxgkJoj1z4lAV98TCTApCi8AQW5YEwnYcaTd4QkAqYZZBZVA/Y85SnjQciFCko/hZS3RJEi+Mf7F6KA1Dz+Xnllit9iovcZFZ4hNY9Jfb2ACsxbSgRfT4DAvi1EBwQOzLXGUrAIpx0HTVBDTIwQQZRcTvwPQ0RAm/3D9+UQLiQBTdwSTjBc5kUQCjod+aUAC5YfMFjCDGDEFLRC6kGHH2CBNBCEKuRfo/XEigzMwBhdcgRAYjUTEFjgVlBST8RXT2z/WewR4IP9X1Qk4KERROqpXIH9Rm8knm+onUtwSAOBV0twYE3YwzswoUyIIU2cIEm0oBu24BA4G6CoAa6k1XMsBBOqwnoZx40thCnIQf88ChAKYUMgT3Ic4T9gCqbEisrRROwRjkbsHlbogGpE05G1xB0wgQwwQRmUweIxACE2hAY2RASMIk34g2s8nBqqhsRxH8GABEj0UgZIEC3OYgumjBrMACXsQwuUXBhEA4OkAh4cBR41n6k84oxBE02wQLg0YkddIUn8EY8N0qrhhMJ0m6nEwhMwASfKQBnEAhGIFAMwgB1FwVGEH09UwELoTEoIgzo2xAcah9QlB0I1xCze/6MEdQsLGgKgjMUscIFITYAfeAIcMIguCAAIDIAsvMIr4FEORc+M2F10FAEjqhwbuMCKtFNDSOPcEQSCOcoJaSRNtJCQNYSMJMcZEAQTXAA3lgAMJAIXzAIzpBUoTkApRYEKBIIKbAPJeEw8hpcs/kMvxeI/dAsvZcBB3aPHtcU+zMIscICh+UEdwEE9NEAcBIAFHMIhSEAuQGQOgdtvyBGLVGRPFIEFHF9DKJIU/sNwcKFL/J1LDF9I6CRB5MJOOCNDZCFbpcQOJOAF/OVfMgELhOMs8EJ4UAIvWAIL6KROHoI24AxNOAMZ+gZUKcIn+MonxMQnZOY/GMGM+EUWEP9EUP5DaB6UaSLlUWaA/VCCNnDATDIAF3CBHygBHNBCIFRBXUyBWrDALMxDRxljTYglvRiib+xfVKBlTKylo/RdSuDkQmBIKBIENZGEwtyLIQXeP2zVb+xBLlwAJQTmS8bkPvCBRpTBDHjZdOVCYvJBFaxCDnFmQ5DCQvTCP5ACKfSCfG5mdITmTKDmaSYlQvACL4QFH/ABM0JEDqiFgtKhGrAAF8iCKIhlHjREobBC9VSKIbGIbF0iTvCW9TDnQkhidEAhSfwVQURZn9TECbGdAc4ER0LF93jMIowjERCEAOxRJOxRyB2XcTDBE5RACSTCP7KBNlhELMzA5fwDL+z/Qyu0Ah84qXqMwgu9wzRsgiJ4phGAQTe8RgyYga905j98Qje0EsQ5Cn8yRBYcQRasKZvyUieopyU86T+0wgyUAJJGhBUo6AzwAiXkAjT45kKIpb5FxR6AjG/UnzOySjqRqP4RBKftgIgKV3SSRCYh42/EaErkGkmwH0msiCn8naoIwI3qqBc8gBdMwlYFADfBpff0BAx0AGyO46RtQxwawj5QQoE2KZgRxIS2hCnihD8AW0OgIod8wzc4gyIsxCcIy6Y8AjZAVWcawSeYwQJgQ0+QQEycaUqwaZpmgTxkwT50AsjYWpM6aYEGwwz4hxsy0Sr8i8vVJUFIjAXsAL2S/4TBVSdDfKSlCsU/YEI1ROqjOAfbtd1Y9d+6QIXM8cTDjMQ/9F9NMUQJqY0xfGRK9IbyGUe//EPG1kS9YgUAiGqqCEDIecH6zUAuxMIuBMI2QIMCtKwCFF/xNcQbHEUDLkQixCpAcsE2MAMzJIKX0akh8II8tMTD/YMzOAoq/oMrYoOxWmvS/oOLcB82+IO1MkTVpsZBbes/dFJDpOkRiME/bIMlqOc+GEIngFkK7MM/yANqMhETZcEqpANBvOsW/sO80uu8HsUOKAMjmsLAfsdvAOyMgOi4zYSHlAESRkd+GaeNEgTjKlq9VcoMjUAkNRenQkVyxQTFJoeoCgAmPP+AMpTDDLQCgagFH/ACM3DCKqxCyyaAAoTCHXzsx74BMlnAE1xAAVxAJeiuDPBBB/iBH7QA8HIBMxhCrqarJexDPcqEFBgtwQTr0y6Ei7yGtboiiwzt1m4tPyzE9hIEMvyDGBwBP2SB7aQAP/BDJ4kB2IavmqppFhRCHryCLDhAX9HvP0BD7v6lBNztDhhTRjDDIcTCVRgcG9jhvSxCpYWE2KyQYZHE5nKUcv6DI6VaxiTH5c6EXLWGJIYHTqhNNbyBiAqABWgBEADBFDwBJeQpgyroEiApTG5DLOyAyALALgBANWTEE3SnDstALLQArfKDNvBCK3RCk6YrJfRSIfT/krbGxNH+qqnMEkO44ipGBzKALfj+QxtYcRa3gfiCRCcYAD9AgPiKATJ87REgAz+AggnEQxeIAv06QCm0sQO4gAxs4xMsgQqowenuQyLA6VGQiPJgiAGbSgSDz8NChdcgwNuZKA5NcEsUGUkkYEhY01/GQpUl573IHVQIwJHkgAk/QAnkQjD0BZ5w1hwCCiqPbitQQiUI6D6g3pIKqIAiJi1Tgri2QtCyLU3QJ4tAsW84MU0wQkp0EvoyRBaTxPe2wRZnQQoYQi6kwCqcbxivwhUYQyysgigw5CvEgwm8QgK8whxsQAvwIp+OrSUkbxCbBEGsHkM4WGsUXg90jamE/xpezgSERDKATQq+1o27eDImAEAV9FLmKc1o0mIK8EIG8IIBKLQlJOY5n3NiJiaeMAM/iAH21rPHcO1MtAEE/ENHh0Qb8EMWv7JD54IlUIIt2zIRE7HxGi8u48nmfS8JgEInkQWf8gIXtGhdScokjeOkSLJpcVOGaiHhhoSJekxRu8QuxBxBXE8pQYB6LO9C8OcSx8RHf+/3krEBYTRUWLFxfG9HiwE/bAPYdm9odhL2hvERQJs4dAszeMuSwhRMYOA/PPBM1G/mugQCZDBXywTnqAY7u0Q1Hl1MBM5fXbAD5DX4sAAMxIrghq16LARSimZkhwS2tgQJdHQb/MY7Nv9vX89EMnf0R+fEZXvSQkDA9542Fq8vQaiv+rYBMsC2Mic0F7CARigKXedEILkxTvwVX7NXSOwCCCDIG4CAXQ8SDgyAIl2caZUcAlRhDtUoVNyzC3gAQYTCKuTBNiDUUQrlQmy2R7snQYz2Z5PiQkwm+JD3TKg3TnRSbCMDasP2EWyDOHykJ/zDUcOmiRrsIMXzGQ02UxQhWRVQAYXEHj7K2x0CPefQPuNEGzXEM+BAehjlt2o0QZT2QmA4VFz0P/RqajjD0fpGiEfFJhDbd+cQeEMAR3N0GPODMQAAHjBuSwz2fTOYYL9LcuyCgJf33RGSTMANHgB4PBPExeLE6qX/EEHErL/QxI4wBW4sxAWnxAccNUkEAEtlAyD4AgZswzYUQpqKAQSEOQSQgIZneEOQt4WHxBF87Uy8Y09wHU4c7WR6NlaAwj+INHiTNk3YuVWLOTLANwk8g8YsNVTswhvsQg8UeUwQtws9OVMseGo4+owsNaEfeCCUkm9MD078RCQ0eUjQcxQQempohKgbNUHwHEHgngSnrDjsw+pmNgRcAZlnNq2PuSdp9j+kdvg2RJoThIULQdGmRLD7hiskEE0ULRK810z0amqTd5lfOE7w+ULYuZ3P+piP+SrQQSEYQ5HYKAXnhF1xcGoEtn69XyjQBHOrhoSFBJI7EnKs14EP/zlPHIZqZKinN4QFJNYupKSjSzpT/BWVh8TgLQQACFrDEgSiyIEc4AAn5MEc0AEo5AEJrAIEUHMVl/FCdBJ/HkFkF8I2XMHmkcH7dQMw/8PDlbyjDMJCMIIwT6iHMwR5gwKG53lNlLa0EwS1/wOfzzTPy7zE50EexEMCiAOkk8R63YB0twRyVI9pLTUh3EbS8zhDMD1BpOQ/3LtM9AA9Mz0K8BBJEACO88Q9E8RQI3xLkA8WpIbVk8RfuxtGNcS7EwQNhAEhEIDd3z0BnEHX04Av7MIl7MIuYMAN2AAFrEASCEMzUJ3EnYMzVMDRNm8FCMMKsINqzF5MwMI/YD5BaP9+S7gCyMeERr+3io9+mI/3aGMrmZv2ZVd7z7c+KLx+xMP+z9NBPMwfQxQ1JKeEL1B97kdFjdbo2J87TagKHlB6Q9w3+IB9u+GIyclE9VDiJRhSk4cQqsXEZ3i9TEChdRPO7hNEqRc9U2A9QVjDJdQBQWAABTz9B1CA3u+CL7z/++sABQyBCOBAEiCBHjSvM5zDPwCElH8DB64geBBhQoSDFDYcmGTgOXo1DMJqyPDflW1HjohJ6PEfMmQQkP2DQEfkqjwQVrF0SQICTJkkaNIEReLmTZp5atJkRIIOnTwKRGR0eNThh4NKCPpC+hRqVKlTEwaiehDDPyxXCQL65zX/DpyEaxok9JbQK9eBJ6Ke+XdGHEEP/xBgjVoMKVuoAf7xHfiCIAq1CCMdvGZNSR1PBwn9Y+r4GQFxhTituqJglYjM/Vyt03MOtB56CV0RxAj19MB1oH8MdAa1wlEFVzgeGdiGYJuSA3eH/EdiVaBdwwUEOlNFHAJOCkDRaf7cedCg8YKuWrUt7vCBu/5RgAriqV+Fz5ACnnoJ6uLvU5UeRD/4aRiCguA3XCPNobQ0CgvXgp+1Ie8c2qo+gsYo8CpdBgIEr4PSosqX9wgisLvPKogtkyQqGM2VFTQURrQaUitoBXr0aOac1w5qhiAWkXpNxYOcOaeZdQzCATNkjkBG/4w2ekQGNwhwC9Kkg+gQxxdfUBjuEl92UQKEM15QAgW3UBCvsYGyJEjCf6o46gb1/gHvoMIKK1A+rpQAcKobCDKPKwoRnJOqsrii5R8n/xEMIb3o5OrMfwKdqsE/0WpElYHiOKoOqcKhwJUbVkBCmBVc0ZDFc14kCMajYksoxYhU/LQhKZIYhCIMBAukkBxFaqMNIWWFgFaZYhoJlEJ2ESAAX2gIBAUqhf2HhjwfIyhNgvzz7x8MSkvITYfwygYhPuMkCIeBoh2I2Vqc8oXZf5LV6h/6Dsr2qHCdWhYqRKByS4eDCLABWkMRjMahYgcqVt/BGp2TlkasUQvPbPB0F/8qg6h6MKFr/kk00X9SaSjecpuglzNhPo3RoXWu4pjTkF0TGaF1XOmmghoo0FeQf/+5BQeVQGHkCstqjQlnEq4gAdc8qhjjyYFQGAMFfQMhZ6B/kT6oFv+c4opaPA/yEyEhTjCY6XC1JejZgRD+R+pa8BLiIPnGnUrrfwpF9h+kyXFLqooR2vYpgRraAr41ErJDIXz3I0hqgvp9+CAdlCCbbIeObXYgNh1y+Kt/0EEQkVpo8e9re6VCOGKwBwrhioHMyOQfYYQhiNR/Uvd4sNRRfx2qU1eogFJXMkFYCU00EUQTvP9porvfgw8DWCXIwQALCm65hRxylKAy3mLl7lf/k3KVoE8J//CqBRFEtlB4qoClonqgwOGj4cCnDBJwIODlHixiSADHs5Z++Q0wIfIHos/cTf5JXHMIqcc/xHIQd0XgHwhEhCrkd5AGKkQH8kOE/qJCLcJBjisLeN/DzJdAhICPIKTjioL+EYeJqQKDBGEFCbfADjAEsHQxhGHphOGKGgiDdTVwhRmEIAUkAFAQ3yMICAfiMFVIjVoWJJbgiPWLwAFwIPGSWqI6iJTBJcQaA0MKLayBp841xCArqN4/MqeKLx4Eir5rHELsdpDJ/cOCtHjj4hpiRiseBUBqTCAC7YaEGeqNK6qIwT8ggY6JcSVz//AfQU5XxzlRkCAI/zxIGwP4N2kcMg1wAB69/mEGMySkGw+R4VEa2TGFsE51//DYKlV5FNYloUOsM10SLDUIVyChjX5MiB4PcsZ//MJdv4jABMHmy38IZIMIqcFRICFJY0puLSfwk15Q+I9rJEqJVHkjQSqGBB0s4H8IwdsWeOk1BPpSi5AkCMQOcsgT/IItbJEkVB5YN0LOMD8HIaFUWkMQSBzymATp40B+IBAXpeKZUDkFIRc6FVaoU5cOWQMgp0GQaQByIHAAJBzsYAMw/OEfigjpP8BAryTUACJPcZ1q8NmQbpyslARJQjj+YSmFsUWXMY2hXiaHDlX01IyJigHE5KeKtMwzAg38xf9AEmXEZCbkgakYpFoUBNCIPRUqJ6CkVISAhK9tsyHxbAgrTNjOh82TIBPD4BgRJBY4VLSlBFmDWPg2EFZEww4F/EdDCcIDhLBiIM0cSBtf04xT+MODCFmUPhUE2IQ84h96g+w/8DUQbih2IABFiiSnipQBDgSu/6io3u4RDickxAacISIY2ZGPf7DDFqEciE5T2hCPrQB8tX2KbkUZ0wytwAw28CTpVhABx8YGnAOJDS4J4rDLXnZyAE0FDyY2MVak4oH1TMgZ/bjStFIlqopSbAxAFhXNUiW5gT3KZQ+C1kGmAj/SwIV4z+tGSdIOhqEN4D0UMlnQ4oIVkFjofAf/QuCDADYCiG1NA/u514bo4q4H+cZBJuqQyhJknwrBBQ8amNSj1PcoDfhGAxYQ3BAkZJlSkW1CoNALF4r0DyEIQRK6wVuICCMJmaAGQ3R6EBzP1lHJ+AcpevEPEfRjBTXIhBlq4I8GI8RF3y3hX//BClzwbb4KOoVf/bFlvqqQvYNZbENwgYuGpsGxCZEGWo+S4YGwGSGSlAKcEwJYx455IF/eawR4wAMIR8O/UGFFP6N8TDrHNSoVJsgxjqI3/PyjCIj+U2WX8Y9Kw/ACDUnhVEIRCklHQq+S5goLCFKCqfhB1A0Jdaq5kub6cIIgqPiHDxTiACK8INKsDs9RGP0U/yDoOq70WcRcqAKAg8hgCQd5gXaB3WxnP3sqpob2nzrwDwYQxBQHofVAfKCBf3j7H3BqdiP4oxBj99ohXzhIrgdC7oa4e9pSWQRVwkyQHMDH0/GGihaALW2uyCGudUFIMi+cEFDrmyq56AADrn0UcCPlLJJedVTQ3RAJNGRQT6n3Qbyx6Tn9bTCwPgqeE+KGaatAIfBWCx4CaCeEVDbZg0lkQxxgrwlQpdcYvUrEHSILheg80A4Bh7UGsgek+EAUUgF5nRoigEbovEAV11w9oE4QGFBOIUu/isgp3FIFzMnlCK9PzAnCb7EjSBkDqTpSCggHbxi7pSCOyjigkrapTP9crn+Cu1rUPRABSFSLDvmsoR5Ap7UrpD0JcbcAMPHrp7hALWG3wtkprzmBY/Ug0nY8gi5d6zkVC+UJ4QBCZO2Decz620gJPFdWX3mFsJxOnR/Ixacie0kXYEsDGZTtCfJ1gkADPrSfvArwoHWHEEBzsq68CQZS85rDA+EG/ke1B9CQ1W+eINBPNeShLYCMR8X4Bfr7QPrueoT/Hfsz5MMMYtGDHgQi9P9AeRRUEAj70yBJcgD+QeZQIOWz+uagouYIgvn0Tc/+wU2IwPyyjQ1M4f/agU4EziF4D+8ix/zGTgaurtkOLyrGr/zUoto6oAD+gRIGQgmsgiDKQSGq4R//GI3RJuEfjG0SJgET0k4FWCAWUG0D4KPhDKUIPvBPBlDskA8qeC7euO9PArAHL1AhiuAOEgII6YTU/gHZmPAq5sD3/iELD+IJ/qESSPAJSK0cWBAGj6IMp6IMvUD+RgAqRlAGZACffm38DuLR/uHmqs8KD6IC81AhSm9OAvApVDAqPE7SeiDV4JAPp2ILCeILn+AJVCDt8GkSWPAo+OAfpvAf7u1PBk8hcoDdFALVAJEPv+D7DmIJj8LxaO8fRC7fWmoHDQUQRdFe5nAPp0IDB+IMb1HSEJGMEtEh+q8hKoEFpuAf1JAS42oZ1BAhykENvWAEmOAJlkAVD0ICDUUT/5FCFvPQCBNi3pACExAi8QbCHJ6CfeAj21zAAUWtMJaB90iOKtaOYaSCGBstsghiGyVqbRCCF4+iFhECCaVCbz6RKtKvIeLCIYzxDLkC3aTuKI7xH2BwCmYgFwhiBKEND31RizgwKqZxEf7xKbKxQLYtrjCB97pOLcRjQaaC7KSiHxFCI6dNb35tGqMiCv8hAZSPE0wuIQfCITmvBReNKwRR/p4gERCC2HwR2Mgk78LnIH6t2kAy1UQSn+6RTtIiAFASKvYRhjSyItnuKv4PKmBvJutjG2IhEhsiITvPBami0qrBC9qSKyoNLqcABibyFM3PAWquC4DtCXLAArBSLf9ybSWnouGybU6ksiF4kSqpwhEUQixekvJUziQJAjAHwuQIAg4x7yl+gG48bREdkyBoTwHVwtPYwA3O8inQrfOMjQWTsdKO4S0Voi0nodIE0QuEshhx8yi8gBJ7gAvY4B+6ESmHEyFITTjVwjAHY/+4zdkmjuR6bQ5FTdy64h+20fggcyC0sj7Aku24I/64YvIG4hBU4AFUsCQTwiHLUADgzjz/wS0vbScTQhmL8SDO0yFYcAc+QOSOUyqehjj17S6fIkC5Aji/DTHBURcXsz6ccyC+8Sf/ITrzUG9QUx9N7jL/hDsdAvYS4hAwriF4AQZ0Ew2LkQW9gDYJ4jVjs0D/RBQh5hPdVIAXtAHWuO4qyuACofLZLpIJtfNPthGQCNEhShE+cJQr1gA9CPIgnnBO/i9DHYLfyG40/yFK6/FMxCPZVEAFC6/w6mMSVfQgeNPS3PM2U5BOelJLBhQp7M4sEkJHU20W0LTZ4BTRwO1A//PssBND/0HWmvT1GqLahOYoZuAfpsALtrQ+4HPvvrE2f5IZGRItGW0ZJsFRj8LYAMDYfLMbaZQrlFLfuOAfZsHa1MIC4u3mOCA5Jc3kYK8yj6IO/wSQ4uD78FQqgBQqjFTU+JQrqq0AiFAhMGEE+AAIDLXwVJBFeVIhcLMM9w5CAeAYHHQg5hMphFI3p9U9/wliJ3ug+qqRKwZTVkXNU58i0xDtVI/ibDQVn7oSPkoyHhFkXZ2tW+kEV6MiSomgK+HKLwJBBtTgH3Dz0gqv84bVC3ZgCtJO6lTQC24zNnsSNpNxUhOiUgkiQv0OQgdCWS1VPaMAXYKPIACgFt51huqCSB1iLKMi7BRiXKeiQNXCXOEDFeIVKgBh1erhEpSUKgJASP8k/EqoJWcIXRIAKkpWIf6UVyOHL94gFqZAKLW0IS5tClggF3agIViwNasVPQnCTO9TWSl2YvviIKYFEL5WvA6CP+10KoCWILqwPloP24BtZZe0IbhB3RyBICUzsoguxAQFs+wFo9yRIHa2If86tD7Q5TMLRAf0SwDegAVGADcN9SC29AFGYAQMoQTjs3EJYkvHVC1EtPMqbUwx4TaXQRmSVQAidBcOYd4OUCGigGwRjQNP9ikADlT/wXWR4lSXUyrsFiEGt4hq8igwj2/L5HdbKiyaja1sciqmcyBQbfoQohEE4AuMYQSgNiGG9R9QUwVyYSL3FXMTYnPnpByWQSgplCDm0wtQcz73zgKUF4a0lQnRtj4M8Sg88ilGj9U+4EoUQgFakSv89ud0z0HsBYrs5U+BrV2fwgKMQWAH1SEMVQX4gBIsIRi4FxkRovAw13GX0XIVogDK8XFUdyBsVNTMtqU2jmT/YWR1LWX//8F2oSIcY61A6NYhIm3pPFYtAnh165ErGmEXekBxGyLtKFRQgcEQ9LVFURQqGHcqInEekTghVPAsH2A+YVAAeiD3jkJMbhgpUM7VqIJmD+IVU20DUvgpphR/aZIf6SRiDQ+HrVB362MaAMEqpmBL024eM5ggpsASqQAFuQJapWI+t5QN67iJj5VMIXYHPOHQpAIENtRQfJbVvvNdBeOEXdZewnggVngwvq6ND4LfzO4gCu4paFghirIoWyoApI4JCGKAzc+DdcEXjEEFoFaQj0IFqCAXjKEcihUpqmF0YRB0FYJxhVUFI9IQZkCODVUZ6DiQq1c+0TMQlgqLA+iT/56CExVCfjXuAvUXIZAUhgoYIb6wlOOqYZkQ1eoKBWJBep/ih2egmP/hAZhYKgBgEsrhnQfincvTIQRRBQwhgo25ngeCmwki7ZC4DN9g5p4ileUvmh1iYkohlP8BF17gQrHti+kxriAwgNYAEQJatI4CXQko0ZCi2irhC2t1MG4WIchY31qgygjJE3pYaRUYoBNCUNkQn6+CnpVhS8sBj5GWIByPpw9iB2Yggv+hE3qYGFGzE6jAENBAoJm5mSGUFkT4IDx4IFLZRp11oRFCBIYh9QQPouGGTgCXTmgNox1CAZE3d9UCTy+uW0VZ3+C6AKECfr0QIeRgNOWHBmD51/84GiH4wBB8Wi3OcgrUwIH5IJfJlIgJ4lcNYSAMIReQVgXVQF/LwSqoIAWqwKlneSDE9x92Aa6PImRdb1QRwqFZTRcRjQjIOiooGT5QADJhuEAqqxZDW9caQEJAmCCGdiCEwBOmgLOfAp2jYphV4Dt5egSCwRIRe1//eiB4mp0PohMCu45HYJYNMp8PAgAwAQSCdyDwhewSmiq+VexK+xKfAgLbge7yUIxFGikSYJOfAgCebo0RBJBsmyq8m601B6MaAGFKYAlKQNoi5homxw7WgCnkmCr4gA2b250VQonRwLoZm52DIRd4wRjsmbH/IRieoRoMu6md+ksswRJmAGr/LdEqZqATEOJL2LAxF7gayiEKnqlkeTQq6HcqTjuu3PcpHk7USppA/2QRHdnXzJt/KVVi8XtuniIN1uCiHGIOT3hO9lIqaGAKK4EXEsEPeEF9AY4G4oAcVCC4kcKYnzshiFHBpyAW+HkHoDsYHLsKgGEIhluwi3ogAqGpE0ISJHwGqCAYggEFHfsggIGCt/m5q0EZ3i+b6lHnrlHXqrlAthgpvPrhfBwhCEB9r6LqRnCVocLoGgIC61QqgJErJASuV1XU/OIx61vX5hop0CMHSuACOkFfpwByYyEWnoAP3MAYnoANO/kfPNkh2FANHkDB/wGoY4EP5Di50WAGRiAQ/1rBEBwbDapgCL6kIdAADYJBsxEiCLxEEv7BqRMC29uH0A8Ccou9sw/C1ncgClAABZQkEJ4BBdruH8wb0epCCiBLb7Bz9JKzhe3qIMIVKix9Ke1wMHTuCT+6QAxe0owNpQdjD+/Axl/YIf4GKztd17hjIEztAlRgseexjolY2JGiBIg4qAdCBWLhH57B1g8CzqtdzqngZez8HwT9sW+eILA93JtgCKiA5vX8ILLAAMZ9UKd9BBg37ZCbDAGABYnxFwBp6epa1CB9Tnj8TzIdIBOiIkVwq4s0DVAd2qg6taVU166oBXJhsRc7IcLzp/+hMbd0Hi1xULc0nW8h0HceDf+oABjIQBKG4B8+QRx6mMXF/SCqoBCQAQzI4B+GINzLHSH6YCBuoQlSIHtHoBVyoZiD+954cwf2+B9yVioErm0bIunsFLu/Hib1jXfxTiCfzd8GwlNZnrL/ge1t/x9aYZnLLtjhHpgRAnjsvNq/5O/B4IUGYggCYQQElSCMngpk/h/CffKj/yluoX2GYCKDgeYNgMMHwpNzQPkF1c4jGBzk6sjF1hSpQhTyQPXb/yrCTqXtAxCylg/L/ik0EeUivkByYcIB4p/Af2oEqmEyQ8u/KVP+5WgoEMjAGbkgQnR36w8wQ1Wq/JMkqcotgd0E3qoCLJihf2gGCkSDhsq/ISL/B46kaXNgH5cDq4QcmCJFS4g8BQb7N2JgHIENBMLBUzSq1H8cplq9ijWr1q1cu3r9CnYqt7Bdj2FF0YOs2kguj6kY2OGrBbVZW/zLxZOowSkK1fBJ6lJi0o7P/o3s0+QPGZBNRrp0fEvSPyot0VSxHBPYkCGSIBuOrLXbGGz/3IWkQiWDASqdFrrkE9XAM11cJf5LRTe37t1f1/AWyOb3wC66fXMFlHXNNeFeIwUQeAyIhKJEmKv1849XrB1EAQts2PDvg38KHQnMVdid4YH5BMZzKYnMQFuSCgH7dx+YAUmcOzt2OUYTMwFzH1bOOLPAM+L4JE9U5rkUhEAGWBLI/xu+DGTcVEvYNpZLVZnilQa/MWCdVVXxZIJAKVqVYVeY6BaXWqm8UOJx/6RVY1bP5cgcEYnwhBdPgRjSyVEDgRdLYXTdwuRIju3E0yju2CBgV+wsdh9/MlFhCHgjtPJPhP+kAMwI1QDwRiC/+NaUQJeMx9N0UBXFyUAg8ijVIgjgKRAkVjng0hxStcjVFzDShds/S0jlDU9wSDWAVI0ItIxLj/KEXG4n7GYbn1xNwJMfYEI0wgiGDPGPL7G8pYIhhlAxA08PjGAMCr6U5I58Wy0wShPd9OFOH7+OItoYAvEwkC606coVMqg65tE/wTS0A5H/rCZtLMHEigYv4hjrUv8tyvzTKU9LefjPIv/cmZUPInra1bu5CUpXGlLtAa91HURqFZxRZTidVewWVUO+BhfFABdD5JKLSq92YoklBZZmzEKuXnYUXy4VBk4MEYzC1RoxbLLAAjHEoCxPutghEC5f8fDHHyFUOdOW0wYSTBBopCAQFUHI1JIlfOygBDrhRpSDVidipcE4AvmgFhfWQa1WKbp9oINLAgi0Q1bDHPBPOwdztW9U9QzkSKU8ZZjpVsQJBI8IuU06NlctgEriP1xwss0QvPAsEOD/xOBOFTjnQhmsSamhUDn/BALOVahKxbIucOCiCyv/uCwQbXSF0I16/1QhVIQjTNESFffJFGb/mClYskM1k1iAwrn/FPMViHVGZcEdAjktkLx0zaKbBhqIXTdPKERlKE+V8CSo8AZ/0ShW2GG1DJyXEpp8UQB8VUa+DID6DwbPBALeP625VEUweFESRCeGqEGUCsYYC47nA9nrlf4u6e8/ntChKMiKAcsE4hGPoCEYLQmcAfADjAxkgGeGOF01qmEBJfBPKm8R2LqmAoPgCQRs3YvKAajmlQ3kqHpR2cMFivI1qxziH3b5TQ7mYqhLkcU24xLA9r6yohJapQQ4igo8uHIGGQxkD9cbyASIRwhjjKAgSGmNJZDxjxB4ZGIrQQNgFPKPWv2jZFHRnHACaBUepEwJ4YCQ/5iy8I8MjAkYqEFNEI5SjnJMIhA0sBfueGIFgcyJJ3VaxCJ2l7eBSAQaKGSO1IQIrxeGhQhN7KBUuvA2rWxNN0AAo9pcMg1IinIqTLBKFKe4EGPkQkz/IEWVeHafCVEhFugTyAiq0IdfjLIomnOHOCbmElSxLkysRM0IyvGAaqgABWmgRe7sFBUYaANqJKTLI5e2y9/QjTk1/FMJx/UPHf6De1JJmnDiEIAdYUop2RCIKqbCgvCFjwVSCWJYsPnEf2DhGVN8Cx+GKSYIfGQID0wBqgh6un+oIBBVEF02/8EDzdHMJQ2SipjQEL9jyi4QKAjAixi1QZfoLl1SYeTvcv/zyIcyZ5s8CV9U8qAbQP1DptkUJyQ32T1dToV4AwnDM4yhhodEhZVY3MzkmjCGKhgjEDsYQS7+wxPOZQWAmjNjWAxoh1/8knWpGQIwXSKTIPyMMhXcwSSOYYEelCsiKnUJv9rKG3C65Ee8sZrVaArXfwRsK/aUCqg+EBU4tK0oZhmIJYVIIuLxqw5niAUVpzJMgWTgCMkCxxgCUZgm/OKAanEZ5v6xhXF6JXLIAodpJkOFIahmIGJiJU/G6sUd6FEFLDDnQ4XBo3a0Q3qjBKdLo2I1rhyWJ6XAazYb0bytyNQBr7jKW4sy2IGwUCBFmMvYnmAV8tUhEIQYbmSjIo7/yQhkAQMBBzh4gF40fiVzZOEcLuywgCZI4j6rfeBQJTSQOhLpmA8ohxpKYAUwinINa4gGj3yAPDxFgCwlwFMmVWqoECr3wXTB6UDMIler0BMrKTKBcbWCL2y6hAaEKJVAWOla+wbBvgKRzEAwZ9XfHNCqUr2KHd4bhiFkgUzizUoQCuSzmBgiGLL1whRqqxABi7YowdFNm/LaG6nE4A50/UeMoCxKawxkecqVyp4EMj4sb+VExMubElJRYlQK5D4oxtZAvpov9fIkxgIB13db17OisJKOP9NZBafgBS88oARCFXM2E7xkqVzZ0LlJZG4GORBnToXCUQEVITBkFQtj/yVDL9gwX8MygapgMw4/BYyYVIzn7tl0c1GRKuakyjPX3vm1Jz6xWONHmRmUwwuTKEep/DUVTgwsXkUhJ6NdMgxPpZQrbrBKcIPbFWksuQ50AUFWlDiQIrikrwN5hECW7RJpd+WTVnnyVxJQbLCkQQluqC1sINvjY/9DoAZYcVhWc2vUoKETp+P1JFTwlq01YtXyVumlybLXmA6HLgTvyqIajpUXmqCvXUCAGflFvq18byCa/s2HuSJigYThHyiIBR/UEAvXFiWWjI6BVVQuFWBE6McrvrWf0WAM2U7i3xLoeMGLgqNGhgXRPFIyXTb+G2kbR0nJ47ZATvGPkbtkFv+O7ooygM0VJZpbIKUQxVXYFBVPRyUNNIhFK3IQC7zkxwD60c9A6h3vPHdWpSiOpVj1/Wdee+GGWtndz3VTzRINNyza1naOvA2+gTQY01LB9j8cfxWoFwXcV5kET9bqFYh3pZT/KABWokAJFgDGEmGS+ZC/y+IHwp2Vk5sKbVg249jrhsW5iZDqVhxkykxLjxgEQXRdoq4PdqUULvBKkzdgimFf5QLPK+JWNB+Wg2NlkxsPpEsKAKomY0XbFgCCz4WIbc5jWtwlXIYX/vE9SP9GFOznTSItkItYfGkgwSB962YOTNzDHT/8n2pUDlhjugFzYVFzfeYqMzAF5bBRvhD/UgNBInfCL98gaVMhdHyyeFghBIwHSQCgZNZHeG0lA2AiEFFwLr4hDSwlROpkeLvhdV4nEJTGEyXABJz3PFjhBn/xD6TXGpE1McAQXjwRLXHXFbqALP8gZ0a4FQOYG3ZnCWKFBoawQDtwfgAAAijAPQ8YFsXXFcGhfX+nFSgoFRVTdVZhFis4FS64FW+QV06HJw0oELWgFV7HWyAEFn9BBbywEp3AC9fydgZQBUIQAVIgBUWxAk3wg8LBWaXRPfVWb5aAdwh4QVSICHDBGxfSFSq0O+Q1FcxXgzlSTXMISYWFFaIAbV3hht2DbgunG1gnFd9HLkUBfWjIHCMAMV4U/xWS4IeaYGCgNBDNoAe49Q83wCy/ITg5knp9WHP1xhqd8Bc78ACTAAAo8E5TRyITEHxFkYoDoVvuMg9s0GwpRBVdKBUXIEn4UiOB93fEUYr904tqEQuQV3AA8HtTYTsDAYrW0QqWYAhWABspsIctxnYUsGCsdhXAGAIhABZbYANSgQN8cowPlIx3xyVoEAiyMwmYcAa1QG0TkHE8YQeWGBViU4GXOBBNhBXm6IW6gXRs4Seo4BJdt44CAY8sEhU8tRU0MljzmC+2VRRA8BYSAAQSsRxRgXRXMZLCEQv/EAuU0AqLsj4uwXbiIAj/0BTv8A/noBUTxRVgUBJXcYh0Qf97qeYS+pGMQYYGMxAIOzcJIGABxlBlAkE+g5gV9ygcM/kbRxkWVcYWU+GBXlGP/wAJBOB3wnEiIRcVmyIQYKJE7aQV2IUni+ISzWMbCYdlUSAQMzADVkCLKfBAwCA4koAE72AP/1ABWmELObKQYlkiqmcArdmaPtMJlKFRO6cCuTBD2NGRu3QGklQU0JAbCmAdnjBd/+CKX1GcLzkVjlkjTyADL+Q7WyEDdskb4lcUMDAdPPkv/yCK/3CBUQE81mFddzEQ87dyFOAM7+APZHGau7ECu3GMRZF6rumawBCbMHFMO/cAT9AB3fQPoEIAV+E0RJcbWUNK8uYJUlGUR3f/MItgmOMoEDAwSICwC5AUPtZnbQOhEJgXFazoEt/5D3R5FR8iFdY1AoeQlEjxbkURAj/QDFcBCwIRDUjAFQgpFXpwFXCGJ/LZmk64QCMwCYEmA4nwjyaZI1/2D1roFbxZImAji17xnNaxnTwxhk36D9RZpWShfgNhpTyhhmFxRF1hbL/lEksAmWYIXf9AbsKxpVRhSkHyDzNgfxJiAOKQCS1KDzxxpy5xNl9hCzRqFXqAlf/QngcTXjrKiPo2Aw8QaDugAjQAh2NTfNrAFS/UiWNjbPASpV6hnJIkYTXSNVuToMmzpQXQqTSSPOETI8o3EKb6OAyTA5hpCf/oEpkg/xCDyhxa+Q+IVxSucBXvyRucaaj1Fj9dUg2KygK84Ad+EBdE+g8XKhxIeqRrcxU12FzWgY7ZKWYf9xvfs5cCkaIDoQxv8FEGc6n/IKaK53xSEQDnlxXjgJfJEhVxMYa88w9RkAuj5xJXAKZRETlgEQ2IJ6NFmKOBAxSsaagEklGA5l9COgDYwazW4QLQuhW82Z1akYgqZBX3aCiR8CgDmZJcwQYcII6bqBYrWKnWwQIZ5nm74aFY8QKLUrFbAQK7QAB/EStkgXjNIAwRkCge+xXQZxU9qBU8U4w8wZlHK5+80IiOpYBAQAn8CRYPmxUYezBU6xXJlTyWp51OwSPqEv8cg4kVjrmmW7FowsGbrMoc43CtibYbvlAFqBJeLqdTXbGnAtEMuIEsidI9ODoVRUuw14K0rkkFlsBv/fUAubCHZYsV8wBJclM3xykQWyO5baWkV6GqfEIvAqGtV/ENX8EClOkVLSutMegSY7uqRYEBwpGeXaG3WeFyXMFjfOi3XmEASAusBNIJCFgOyvAEsupsUiGgWlF8GCuxXyG6PAG5XtGlmsSXPJGbW9GiDPYPaBsVbHC5XbG8PAG1Yhal3LB14CNPTFAAlKcVCya3X/EILgN1MvoPbbQbuip5V2GrfDh7tlu7ZImADIG4/9BEd6A5DdC6PIEPH5ob1ysc22v/QgTMI4sCmVsrtVGRqTXCoAJxjR9rHR2yG+e6FT4LFriQvpsjl8fSr/nqFfVglVixurohOIATFPZ7tHc0BfSDuC1wPZFCfgNBpbqxAcEhB54CIlbLE2CztsLRwC7RAUBsgdObFYtgk7nRkTX0llEBgyWktWrhO2VQAmLqu1ehUyF8FQIbVXxSt/BCtGMyJi1cu0FRu5bQCjE8BZTACy3QTQc6ToCAB9rWpFBzPGDhdzxMFgcQvDwxQwKxAUg8ECQ0xDyRrloRnoriyBF8FcoAySWiuFsxeGKmk1wBojzhO0yQxSUAyk5kFU7gpzwBxv/AwVPxCCfME6nsFUW4CQIR/0rCUcZ/GxUG1cJo7I9trAZq8LSPlKx1EA0NsAZxgAfOKhxsUHwjey8DsTQisslRIZ32aMHWoQxdoxWVKxCD18S78SIvkr1eQcdkcbxFsSkywARl4MlY/A8DQCIVrKLlKxWnTJDG4Q8BTBaty8q5UbSzOxBD0MIAncucuY9qsAS8wAuPFBfC3AANYMyGIgsfmsj5Iqlf8VzAKxCBnBvY7BXVCklssMVTcbJdQyPUyxzapoZdGrNF0ZFx4TsYPHzUfBXNls5lYNMlsIdhFhU04gHM8rouoYnoOxCDyMEp7BVGnavMcVBRIUeoMkEA/dQpMEEVNAIzIMc85QcDUAdrQP/McXAJzdN+yRMklDAQVDMO0Vy8RSE2Gt09DTk2IZsuYLsVnRLO2ZRxZQuGU3EDYTGDNY3F+8KRjlZEFiAOTjAKzuAVP103mlAUtCocTR1HMxFHUk3ZEzRBQcFvI3AB+5DQHLkvDF3Ml4AHA/AKoaANwwDNvHHDIdIVyxySLtEO77pDYdF6BsMJch1x4mm6JYLAWWHAfPIEFzCDNs0CRBBqs9DNAhEI9vMPP4iYf4cLSdCV1iFHLmHZElTZKcBvM0AJ+8AF4zM+A/AC09AA05AGAfAGXMABbnAI6cC4Y3OyNcLWZIF0LFDEjAbXXqGhv/G8TvwVNDAQr+DRW/EETPD/BDYtAcbNDAj93eNzoBbwAhagAgTgBLEML/jsEjyA4VEhoz8dgFExjHSRAaqlWtkdBDPQCi2gDVRHdQMg3uTdAGkgACqwKmi3CvMg28YXFiQUzVix1hmd41oRqngSfAgAz68ok3ysG2/RyFaRIlNcQuyasVIxrgIR3Ewg3EyQA8atDYkQC7GQ0NuwHRYQBQtlDHOwDYmNygPh2K4rFWPQByHwB+vJE2AgEOzwCaRQFEbwCVjhUFxR3ZINOBJE6IWeArBCCbPADLPAAbPABRMwACgAB8XsC2kWVCygDe+d0QXME9mgZU7eNGIz0VpBTdQc5FYxLkPOE/e9fVlRdVPp/xJgBJmgq2zkGxVsSMVY4QAfh7UucQFXzgRL0AFPxAt8QE8jwAdwnAssoAI9kAvisA0UIBAEmi99/gmfoAgD8QdWce1GMDY8o1oSFO6WfejZsQ+L7uhcgKyeIATPsCpTwB1TkAM5wAXVeuq6oc0ZXc6ipLWq/hVBKRBN7kSLECnkcwa7gdtZoRc8wVO/PeD5Msj/0K0DUcV/EpMCMS4rKElZzgKJMAGc/W5JMQN8MAMXkAicHQyo4g7sexVBLRyf4O080efe3ucC0e3WUdtFAUeSlQFZ0PM/v2OGwAcJre6czQuU8ASLM0X0M0WlMgvVGrx/+Q/q5BUvMs0yXQpGSv9sXtE13hEVVY5+vAHwWTEAsC4VrB4Vd5LfHG0V+f4by2odJDLI6dQIbEH1U5G5A+G4ETeDJdACXODoeAEbmPkPfJB2LdAKJF/RJWTndk4Kej4QM08KvfAPipDtJSI4gT45cOTznQ/0vNAJrQD6If8PmqmZvYz6Ta8CXJAO/3DxGigQIJkVSzGhzJHWdFEAgGUw+80T/GL2Xvg22SgQt8m/NSIA6RQJkZDXv0GOT8ACHcAFXMAGzGAIsYCZ17+/KM4HhqCvntIN61AUdvAN3xADihDzn1ASdhACMD8QZuAMiZgbIy4VO2/dnZ8FnQ/6naDdAhE+ADFjxAwrIwqqQTj/MJixDbKG/YMYUeLEiJgoXpS4A+NGjhg3dIToAOQ/PyP/fQHwxSTIIisjCsIIxGVEDhAtgLwws+OriwU6TPgHVKfJDi0DBIiUNIAAL14u3lhp8WKJfyxydOCSddU+XjMget1HqRWfscGAMQoxZqSzobg44vIHsdunPxCNOPsm95NdI58+jcEG1+3QjhmyQBwi8XCWIVkMN+bVqVWKTnxmWLY8YwlBgyNG5OIFLNcqWaIo7vkng6PGji0lutYplfBsjCojCqAtUcK/F/9uXgQ6gAHFRv9wX2R90ZQpwgUiJs9tgmLJjRZld2ROkRdEAQKORgoAoKmXSeT/NVICMdQ//1QYr2O88GRJh1kMuLCBpo2XpVjBLHUdq5VWDBiCBI4iaAuiR0bC5Zsf/jDCLluweSevezb5J0K7wAjhm3dyiyiFkRbLosQSM9gmsk72yaWVGVy0zEWBXvwvBRsReCUeiDSASAGIKvlHhec2ym4iIf+B7p9YZqrmnyZBBClJiExhIyLYoIyJo0WgHI6TRdjYcqUCcsKyTJeKRJK77wIorykVVJhEgEZeQIA92vZ4gon5ZsmKAQZC2YarfSyJ8cUgMsjgHzo6QnCmBRfECJtHcHGrgW4kUqQbXCCFyBkzFDECDEUAw6bMxDhKVLESj0AxBSpa4YWSysbCbAZDLLEx1/8UMlhFlC4wquQJFYoA4Q0kd0D2nymCgijMj/5JBLmZoIHoPTOHhIg6idioaSWqlnCpN5egwmgZifAgkrkwuchoIyZSUw1EkSCCZ6Unjf1tpG6rDPIfAADobqk2p2iFEj52iUQJBEJBRYH2/kkAImo3IjMi+ehjoL4JGNiGH2Yy4IMPJlykhIsjJJJkokb/YetaidziYYwQurHFlhi+KfXDf+6JIZxwJIXIrcFyS3WiwxQ7Qp5/ski66QwsWVHWVgzhIxdcIUJ01xSGSIGfPOL5lSIZnvhnhC9AQDbtJLMLs0xO/lGmWpcvGmGiDZgb7h8QXJpEJ3FNSuOfADoCAKP/tmci+wmysZy3oxYgKvwfTADQaHGInqh4om4lks07AcqbZArLJMjFGGO4CEUbBVZHJQEFEoDGjcIF+PcNZVQowbl/coqPBYw3niArZngJGbPJTGpZirkV/AfSR75ZQ+fmI6pwsAXd4nRoLBeTSJ5tlj6CaXlYNYAPXjJI4Xx55EnVMccyGAL+VV7x9SKymRjhDbWTTfOffSN625EoAoOO8Ggi1pIIlUBSCo5YADpv20hybEMRFiyPIoEjzHAWcTiK7MCBFMnFtRpHGD5MBDUz6U53jqGMSSiDBbEQ0gjMpw1OMMxhq0uAC2KRwn9hAhMqkMGYxnSB3vlhFhzISlZm/0G8WhnifBkoBEhaZsGLYO8fQ3NLXCTij6GdQntlOtk/lHYyMv7jCGcUA/uoQAVe8GMbSYsIiQxjGGS8wgGiGKEsqoS5J4wAE/tDVi4ScYd/DKdIi9jcbBhoEg54iQ0QlIgPDBjBmewtIvmCkgAJ0zeK4CZyEMnbP0xRk1AaS25JasU/LEdFjBwHJfZziSlTKABMAOEB5fjMEkagBiuo4UVc2EYooLEKBcyBE3fgIQDe8EMZ5AJzF8DTE1jQAxVQcwQsWGKtLmMAxKwlIs5QXqf+Ec65PSoiWcTFh7jIykQpTWkQ+R5FjiCGM/LiVv/gx8nEsM8zyqNE7IPA1/5Riv87dgGPsuBEAZhwAT6MoAg70B+yRsALLoTQfxCB5D8KgEmXjGM2ifzHJCeJESmxkoK8MdwAKKKDlXxyIovI6NzaFkqTgqQmQHlD5FKojCk4gqe5IIgadjlUK7QiEfvQhjF7kMxq/JAFmHMmEZ8Agw7wgheJyApQaTUDNDxxI6CYCFvI+U0LWlEiHwLa0CClRYwsAErzjIgY/iFXMyJjnvJIgSHEiIzv8ZOeZ9xGHfPggDsS1qBdcEBC+cgCIExhB3WLlVXrdtEwjZIDq1wJjwwYNo7UKSL8ogiPFlnToYAAXRthQJ1UGhEadFIikZhb5hjJQSrK9h8f0CBt/bVbiCj/QwsP+G0sKiEQFw1VqAVZQixAk4tYBMIC1ahG6FgQ1VZcoBWxYEELmKENLvCiFZIpy/EQRdqzziZn/wjMRlxBxTByZJ78kAcvqGCIffAjn38txBlXgYw52BGxiIWHAxC7iCeUoMAskAAlrBrCXHChBxBhV0xvSxuPSsRYT4KIHF5K3uVx9B9nGEkcNlKckSCAphspIWE2RxUOg8SSE8kBEGzpCAFNlBcGQMMMpkBUgsyABSFLBC9awIt9DGEfR57FPpJsVatSQlZikUwnttORLLzTZevk1EjiwtZzRoQHEllADMAIkfZSpA1iQEZEztyGIwzBEGy0bxvsewRkrGII/7FQgIDtuOcuvOIVHMhFJbbDFUoYwhCg4cKS/kHIf3CQXS2GdKQvgkGMAOI8gtvI5nJRUomkUiIq4DRFTryRiK2GMJ6NyKNBYK0caEELtlSBJczyjxRw0wDAQEMwZjCjy7yoYJSwhIKFHVlhO1lWnTC0JcaLNUljo1QreQcuSvVsSZvxImlO81znigw0P60T/1HakbciDl7MzwSrAMUcFDDMbQwvVgbrhNV4IQ/71m0Hy+LCLCRs0ilH2pTVJgxsO2JRaYEI1Rzpwhw2oprj7BYI8ZrIg6NEEQHKeBKB4MUQeCGiixjAAPM1BLI78W1g/wfYwg72u0ueqO9ZGeASmf/iyyVS5o3Ila7/aINEIAARfiADryeH2pMpkYt4T40sxSuLctVnRhJAIAXA0HgGeNFuTsyCg5acoMuGw4CaLGK1rARBb27yt5MuDwcXcencIK7KEkdkOB9YHgzWHpEXcwSBEJkCEJZBOS445iIi4ngG2OfG9bGqu+lD/MaJTG9+zPXmMl/JYKQ3m5hvhOYUsXlccQ4Bfux8Io1HBjLyybVcDN0SpR+50Q3RHz4AW/CNl2sbICCPXFCh9PJmhr4fHREYeNhl7AqlUCA/fBG33Q0gSTHbQXJwkDhAOiDBTcNbsnbbbsSS/67KP3IQJGVgQgCEMGPRdAKBnZf/H6ugCDL/cj58iGwBIuvViQ2q3ficy/4fnsdItvEpZ74yJvHpQ5R3yoJtUBoxsD9goIJ/+A9esBp9KySKiAWsM6nUYj9WYr65yTp3gRKFq0CK2L64CQAsgIgr2AaO66aLaC/807mJQAYVhIjDEL+ZWJkOtCADxJI0Wz98wjYyg4ibk6sj2JohYAYxsK9BkbqSGLWZmBeREAmeWIkknAmVyEAahAiVogCOGJx/gAMoUQnfE6Hng7wKyoHtmwgPWI+JiB+OyDkXNDOcMxoqpMHH+4dsM785HAr8y8E026eJiD1+aIMWNEB5EIcUyAUYmIAJuMDZMI2VCI6O+DqQOC0qJJeVsLSN/yCCf3hEikAXlTCWHSAkyyGg5RM+kABDDpvCiQACBBKBf4in2TAQA3FD2cvBF8yNyoNDKJnFHFxDnYBF/ZuI+pMIIvRDP5SzjPuA39gYjEg7hBshlxjF2SicUxw+ldKwamO0fzg+SWs4LCE7itiNf7iSiHCBUFiF90EfZnMJz2PDaxmrWwQRX6SiPMS5eUIzPwy98LkzlYiCVHMZEXRGk7CISIQIKbzFavyHS/yHE1geldgFM3nG3IAtgXu5LQkFBfA7+JGIKJKzNsi5K4gIj3THf3ArGpQ/ePxFN4SIHFzHlYDFjTgz0ZMzfigEBAiEuwvJivgHgbzJf5jEmdjClf+IRJ2kDZXKRIiUuS0JE05AAE7YhsQ4xyyIIjmcjRgMSbYYSTMRgpHYxfJryZYkjKZbwT/kSLEUAwgYgkD4B2PZBU+APHFYCXF4MOzbiKKUiIa8yS2EgzQInOLjCFP6AruUiFCEiGscChmIFoiImHrpEYiAO4nYG4nEiB64gyj4GzkwSEwsE1QTgF0Qh21oSvdhmvYyyYtYyY5wOTKYiKvsQNUcisYjLfRzwZ1TP/UbxlVYhSo4DqFURogAzIlASIyIAt0EkWWciGzkiLo7KapQAbl8Ob68iH2MCOKUCMJ0CYmDCBeQiFIDkQr6jbC7CLckjN+cCF8ojkYYg870zAz/OKM/JD+wvAivpMEmYL8oUjOMqMOOgE+OgEVY3DnZa8HQW4VtQMvhpIg82IgXkE4qQgFFy6Tl6cmJ2EaOgM6JiBw8QJdtnNDZaMx/ICBI8gAAOsN/IAAQATHLnA1NGglAaIRI8IXORAam6bzO27krgEWQ5AipJAxymsF/qLCOwAD5+wf4kwgxs0UxG1LaGIV/AKuNkM2RyM+IeFKdazoIaEHyQwZQqIIsJNAoYFCQ2AV0Ec6ZGNGJ6E2IYEsogQEhidDcEE+QWAOd8IWI8AUwxQNTYoEKcgnwHIkP5YjTEjjIjAix64g2nYgzzb5u/IdE3AgLqIJtID8rpVISoFEI/5BUiFjHnJPDMHK5iFjSjWDNKzQpW4QIJJiN9dO/0qSIKMXPpms6UrBSUNiGHZKI49BSl8AD5DSJOOUwcbhMl1nF2RhTwrgEkxhWiAjTMvERnYCtWo2IBwPMYM1MnVCmQDCGzgSFVWDVSZ1S8pM98nNNVfEnFJwIUqUI5VEe1rwWIN0IUkXXa1HV83MJEpBXZMhWWDUGjcC+6KMIQsUI5oRDPaVBUGUl3AhT63QJTwAxjEjWlVjWizBYiODXxtTVMqnEifgCTLgJtfwHHAimVaADULhWSaXSkVW/MzojqBwfExGjiNiGQoiiZIAIDKEIcoUIlqo21PyHusAI+cQIYP+01I14V4joVLAiWhIABaOVVwhgBI+9girolyj4gjWNCLfsVWPlsKodimJFSH6FkoXlsLzMSZXAVUzbRmZ1mRD1zYkAv5WoO/C7RK4dCgSgS4moWH9JCYkwhgyDCHHAgQEYgiEgQds8P9jUtn9IlW2ok7ODCJ9xh0xwB4hQi+WpgX+ABZ2oXDMAyaMZzTm0USa9v0r1vPxEv4loyaM1XaQ93TxIgHhIgCtY24iYoIg0CTy4hGNdHrSViDrpARTgzZzEjQCIxA3dyZUA23OBiAz9h2JdidaijRDF3Qn7h9cFiUB4gzKlDUStQsUFStbyBAqAOwKQAwIggCrwhF2gAV//8IVL2IVdCAQsoAAycIJ/MIMboIAt2IJNQIJmOIdx+ocKqID+lYjIhbxBCFInKIRNdUkDbEH/vL9HNT9KheB/eEUJTlV5Rd0LBlmQzYOvcR3GRF7ckF2IUF6MGNY43YUAmNjlEdh/qMiN2IWGG5wYPi084N3hJa2EjYgJtd4yIQBCgDsssN2JEEjhvRasbSWJoIE6wABC6GEC+AAKIIQzoGHzVd8AQIEPuIFM4F+W+Ydm6OJ/2F+I2F89SIIViAiZ/QcBBonKnY3J3Qhq+IcoujzMm0OOhABZHFkHhmBWpVQL9mM/Pt1ABlmkpYNCHl0jmdWJ0NIVdkwRRuGcnJvf/yTijUCBiVVe3KhhiDgESMOAf8AA7O2IuiVWigDUkRjh2YDjjgDikcjkWkjeZ8AIf7wNGhbTjRDlixDBD3hiQoBiKa5kX0BhX1hfDMhitvBfjrgUkEjmkXDjiGDjiXDjZ94IAv5Q+py59IMIowUFSNVjPmbVPwZkDEZaC74CUKCDeMgDEbiC54UIAaphs8WIMb2ER7ZhU65LiRjQoSAE6ZXe2XjTBmDlfwCEW7ZaXA1iiQC/sR0+5c1nM4FnWQY/uDsDFFAC3n2GKgiHbVgFdXYCG8AAJPjfc/iBlTCDi5BmkGhmiKCHMJ4IehiJN5qno5GrbLs5/QOFIXiGziSBVf/IY55uOp/GVnkN6kC24GvNYFDIg20QB3FwgjrhUzNh5IMO2FzFElmmCO0FCUsDBOfcCG8QYVeGCL4kMYqoO6mWiEwWUYl4apAYa4KGElA2k2KAiDpQ23/wBQzYhjxYBb1ehSvoaxK8AidwBWGogHPYX7bQg5SWCGoYhMaeiWZehy72Ypi7iP+lXAKeiPWC6R68uW+FiBbkVAo44fUlBHEgxzyYA9T2ZhrF1j42XXPOAzpQgG2ogkDojn9oyA9da4pQCbOuZzMBa0jGEraka4Bl5KHAIK+GCOWm24goDrmOCBwGsWFlXowAP1imiOOWiE4OZZ3o59wQWBSwhpmgBYn/oGuJGNZLqIUAoAEUIIeLrgIC4FscoAYc0OL/dYYKqIGTXgHMlggCNuONqAGX9uKR/gcD/2KTIOOJoAYR2AYxyC87xDYFXsFsmwMyWF/gxQNgXt8zKG2+JQPPZMpC2AYS9AAcwAFxIAAKIADsFmEG7wibdQleHomGXong3ggjlggQ823oldOJOOUyEVIsSYNrGGtbJjHoju4PuxaspiIRtGqQQOvsxgi+FOUjd4kAaMj0QAEU6GSoWAEp0AP9TQKIGHB6oAcAL/MAnwjMXoEB14MKmGyJmPON2FGImGxnOIckmNx+aN0jKAS72qczq2PPrs8rFdDNVN9L4HCKZnK0/0SBAHDlQHiGThbBTiaEMLiI756I894bEECBIKeIKE9eSANYjMBhUaeIJeZu1lqJHe4ImIg0SpOIYmDua0mPjcAAUq9AcrlCgeXLOODqiBAxdGBeHCbhiMhkLBhRV3AFPQDjCliHMa+B/r4IPXDpZ66BGtCDw6ZzinCGOr8Icf8BZ2CLZpACKZhcCgiDK5gDQTdANFNgzrtjN5zR+1sFckDfXWB09kYBUJ9o3tUBfr+EhMWCXf8HLIhi9GZvXo+ISZTxf0iKfxjvjaBrTU/hkZhEq8ZxKMlnVd/0iAB5LJF1jnC/jvhJwthLiIBuV57y2ch1iYDW2Sjliyj5kYh47f/miGG/iJenZInQ9H+ggBvYAmj/hzT/hyTwYpamCC/232aw7CkS95WYIls05n9YAQoQBBQIBATgaTozwLEc2W7N45EFhULYBfT1hVpo70Dgeq5vrX7/hzDAArpPeE1PWPVeiRew2dZiXubG8rmWiOBWcolwcYkY8n+oBUumjTH1+Y6fiDAIetpA9mp709mobpEnr/SAfCgpfIjw+dwI/I24+Y5ognBoAjN480FwhZWec6afiKm/+uVpGS3WhPqlAfZ+hhu4gjy4gtBjz87zz7KH1LMPhAAohvbucpvl3QAY1sil6+j/B7SsBVd2ZRoghwcFiWGteJf4fMWXecIIg/P//gfyp4j1SnyJgGeKkP7MD+jz50mI0P6JYPOIMH+XWIPL54iUXwmAoPVvIMGCBg8iTKjQoLWFC70NFDjwhMOKCQEZTIMQ0T9EHAnWQkiuyb9wTvq5Elbh3D9nBF1afFmwAkGaLAve/JfzYAWYOv+tWFFhBQYaxQbW+RdG3JVVea5cQQZBKoSqVUlUvTIVAqhVz/7tCpTwKMI6SgYeDRnzHw2CvkJKXBt3YMiP/1wRxEvwLMiFggjqWHhDoVqH5NYORDGQRtuCN/QOvIFBoTvElgfCuYxQFeLG/wKTrCglJsa1muj+y0Yrm0LFljUmjHOw4b8InsH94wz4IEphKmU2/yO4s6ZBn8YXnoOZvLjBm0n+JWmW6fNAvkjJicMhQkSeBE9JNA0/lQQy8k3zkCGHYgzCBQSTEkRh9B9ZGpU1lyYI6NfCbI1SSxSSZwnp8BFE/xTWmmbe1NLgP6tpplBgqB0E2UATRmhRAw2sgRBsA62R2T8fYmRXQrgppIQONAh40AoHUXRQJOhYlspCAiWY4UBxcBMhIhj+c01uBP2imDvaUWNGJsL8sw5OOrb002g0BVdQlWvRBNQ/TCaxwl8U/SXIaWFQMFCZFNxggxPbeLDNFdqssgoJcoZ3hQeFfJWQEoLs+Q+ffwlES1omrhUSIP9Z5N4/EBVTC1kKlUkQLf9zFWSdQ5FWSmiGuv0DyYMGubYQpghB4uk/W5xG0F8RNvDPGh2C+I+IC8km0AkCxmhjQZwJIcRBUvDXUYaN0GgNIEJCSaFEA2o2q0WcCptQNiH844QZNjxXEU1ZWnQct4o65NNMA62TxCBJ0LTOixKpeFafWr74IkGIeBNJLQEUE0m+xQRwySUENdZWSL5W+g9fIVlDC0SCyBuTQP9BDPBBSAyE6D8RI3SmltHSVxClqV6qmRLuOgwIswgmNKpBo/3D8qrJ/tPqWh3CIU0askX0UbAG2RgYEkAWRBFFW2xhGbGNNIQslKo0Qksj0C40HcwEWcMRIhTh/A+N//ThBBj/A3WT7dRjV6THi3o4+U8mZqwQI8H/aDLZPzUYRHRbCYfU4FGN/sJYY/9GRN1AbwemCmeqNATyQnmj/E9p+e28UNMWLyR34AQ9PbhBvR40meenVsSabm8bTJAqyB4uMWMA//LoQhEcRPqWY8MKa0WwXWOqqf/oSpCugQFNkKcnI6a0ZTEe5DQtUB+0atFwC4L8WmncjPPWBMWRhi5pEBzO11IPJDaUaVeUk7gxdZkJt8K44goFUugwmg4Ud24QOqWpgtF/gNCCSFtC14Iik2qZr3y1ACkgAXkYyc/cnmcQT11NWIiIQ9YcR5uEIC0/lDsI3UBXEGvkL1D/AFfLKrcQ/2SxJiINqUVgZEeQa6jCRtfj2D98QTyFIAJ2EdAU2WxHEB8uhBtZ041udIEYu2hiEwRRnEKMBzNAZIN/DEyI1Jh4gt7pSFew4YEN2PGPP/zDDAd5jtjIhxAzNkkh3DqIHiK0jnDMbiC++ccgXIEBll0IIfQwiJD4VxA/8idGPJTeQhy4mWjBjlIDQZbQHHJBv7wwNZI03s8WgKHdDWQ6hszNLyRyOscNJIWf0YGigEYjpXEjFdfgIQ8NosRT/IMH/zhFBCLgHoq5ZzQkdBbZELIG6g2EM5DQDStgxiSLVHB6vuNj/g5no8MxD24HwWSEolEzgsChMjYYCBgL0o2CPP+HSetw0jF7WRA0ohEhSQhHEpgkjHUokW51BF/LTvOyOPJxIFvb2i88Eq2s3ZBnBimnQexCzYQ0siA9uh8oK6LED/1xhvAbCB5Bp8mN6GaGpisIHiuKDidmTWcFaeUyO5UQmEjhfOZ0iDR6dBlPDfNX/6DfTH3Fst0Zbkj/iAMWFxKNgZxidxHw1PVsRE1ZOiSaBQFiQUSUGThYMwZmMEM4urnNf3wTOgdR4j+UmM6KfJUgYSUIQQ9SrrOlsSB1vAvFpMckJhIMf9fQ1TP5E1NV3PUfyIuRFGCHrN4x8SC/sBFhE9LTg8gGHbJxoo8sQjGaEoSQBcHiQSdbEJ5u9JD/SMxQBK40EIiu9IcD+WlCjIiQHxBEli5NiHtIOBBI/EBXih2RZUgbyxgMhBsafe3UZOaq38oquAZpQAjA0M1uhlGMYEtI2o65xtDGZAWDMEgFmEQPumXCFSsIji4H8tiZFgQcgNBNfsZ7wtQpNUgmrUhlHXLY8BIEHemtCKEiIFmEuJB3OpKGLqRRTINADRDXy29MYDeQH0hjtP+YhmiZCqVXFSTBO1UILAfCAwPrN8PNcEZKo1QQWZ7iB55ihSoRwsuEREMaCU5wMXWxNcYKbyF4TGbMfAlcgjQgBjZQBLUKoiY40nO5BNmESbC1DiSMU47k0sxYK9KlbHEpW+vI/wQ15qZd6oJ3jQf9qHoHUlgUUVgh9z0IiTNsEVjy4L1aW3NFEQPTtbTZzDGRLM5w8Q8j/jcmkIUunwmiEVxEww6jtRlvYWnoU6SiR6YdCIb/gVpY5nkgYL6zRvyLmYM4WFbFZAWNFdJogR7kxMP9YQM24QRbFOQPYNSu+BRig2T8oxe9YIQiuuGT6or1H3sMH0GSoK6GnVEzUl4BO/IBBpTUILtIqHBCPDvhhJTZzx/+hz/M+d9IQ/sfkU6wEa8X55ggFSGpoEhFfYLaCG9av72LQbgRwgrYCHogJG73ygai0kz3eWqZYfA3CMLsf9jZzsWUjYQfOMuDy1vaBdEeQf9++tTf4nsgdoZZKozYaYX4tgHhUMRBqEo3umV1If0YCCn+UfJ/MCIc3ejGJrIF2WNmq50r0O4cLSOMVoPTIMmgRrLvMpoInJsgP/BsGr7MuziwQtHa/oeE/3uKatN7p1rMEGgNsumAY/vZCI/QpwmS5yqp1CDbS0Uaikn2A2dbIVnfkZrRnu8+2/YRALft3Cd+acsaxB9yR7hGcIZnzDD47jc+SOA/dHE7/DvoOmpVq75hCxv0gSCohg4Z15KJHg+kFwTRPCkYQQpSgAEMIS9nuW7evkzs2pVa5apWHdINRmT+HyIY+QqSQDdXOLsgkIgAXbWdNaSnQeCw0UVm8lw3TFz8+0MFj1DVlz53WS3/swnvutofeFjKOtogsJQGLniZNW5rP813XrSrBI3nsh/E0hQ9SAwCAgAh+QQFCgD/ACwAAAAA9AEZAUAI/wD/CRxIsKDBgwgTKvwH6NHAYgsjSpxIsaLFixgzatzIsaPHjyBDihw58ppAViQJrqHYYOHKlRMjLYyG0EKPF55ItkzZcmfKnwJ1CQxQEOZCBQhzAE2o9J+AkA6WZrz3TwhQo1IV3vkJ4KPQpxlfAAD7QqHPghII1ru4NatKjGs9uunQYWBdgSgIjvlnrAeLET1U/MO0g3A1TNV2CFT2b0ogFVHu5CLCRducOQW/uN3MufM/IJ47wkjr8YGXcgPT7MQKKGNXjKAT0lzj0xtIGDAiMp7oYmCoi3cLDHTj0c+/pgMncVbmxSDqf5PK5YhlUMbIEv/KHLQTmrMHgQw2Lv/qnjES0X9ECvZGiPUg7X9rWwolT7++yGPPLwooBkgAgGoINSeQgCIROIkFh/zTGychYWcfUGdxNMBSUWyGikDmYORNKghJw01CPs0nEFhUCdTeRybJdF5BDpnI2W//ICUVWE/MUNBuCJWj4xQqqEDgQm/8A8B/BP640DIDIamQkgjlEt5PK0XgURccmfIgUL8YVIlbMCqoUGwhxeFed3BglGBnEXL0AEGx5SfQA1PEkgsljQ1Uzm53ClQOJsf8kydJSKKG2pp6DobJoQBgYhAKOIx3yk8TCGTKLFcqtEdBaXK0QaX1nUiQdRQFQNRLnCJ0V6ns/VPmHT24udADOgb/08kIzwlKkTJu4uicn//o2tgI/6iB2hS88romoRKB8AxFTICKKqdlGbTeswu9dlG0Gn1gkacZJdAlS9T+s5JPJ/Rw0IQEIfJIHeYKdusUOfAxhY4G4YgaY7spgy9BhlgCLEFwqsEHsHDuACwV/xjCiyXE/hPLvOWMYMg/CAczxZr5HfsPskK+kaWLnuY2kjjhlmxypyJFYK5IxqHbXQktXPAPH7nMmUsilCQiJx98sECQuwaBBtoUM9hY6EDz/jXvv8GMIPHEaFRBxRD/VEGdI1NMEczE/zRtiCFVCIRGEClIUsUQCA8UdtoFGTJCww8Aq4ZAYPq5Q6tjjfXGDoEE/yIULiKBAMLJnrXELeEXlfhTXikBPU1B0YiJuEATcsGF0UoBLdC/A+WgxtxzE0S0JcYEsoMxVVTRxy1NSIIGFWFLosgfTQjUxz+r3yJJMFsPhMY/ryM8hCS33I5761RXTQUww9vyTwgDhdAH9MAYEsTyGRhgiI0NT9FK03yk/Uwwz4wBxz2ZUjReZ5QOxMY/DHp0AH2JIHQJefBsNO4/gF+0ppIyEdc/0ieRqAgkAZPrCKW4MAHL7YMLvDCa0wyRi0K44x+/uIUx/mGjsBVkblMo3ccMQgeEYOMb/7CDHXigiwV0IwTd6MMoNhGDGIiIf2USyDgk4g8nKKIP4RjC8P8kkQKKUcFijjEEJYJggBQYggq/410wgPEMXezkGytC3JOehUBMGeQEGJFZqRykmASGREUmi9RABuCJDQ6ED5YYCCP+EIIm2EISyQvCPoARjH/IbQpVKF/J7KALdzhhCMAQCBWC8A8mysMAA2HkIhvJuUDoAA7fKEbDCDceKyHAjBXRRSPOAxbO7LA+dbsSOhCSRfswgSCzsBJTujaQRCbSIHgcQga20YQYjCEMTXDHGMbgDg6NZBMbYaENGFEIYEAyA8C45T8gaZAgWPMflkADrcpRjR5IIAdaGIgjMvK4wYGSIxowo7MIl4ZzusUnMHkCRZTgR4FQUyGJZKQ79bn/ketxcASwmkIJlgDOzwgkGwOkCOPcSa1SdkRRqTSIKAaCAykh5JX/ENw/fIERAmaUO+/JoUIssJBSeIRARCnCP1SqUoRQZQ332wyDOFAQVRBkBgbIZisMYABgvC6R9ySINEfCHV3wgDvP8ucMIKaMEkhAAAEAxBoUx1AzfkggeCAIcjiThnZWVSE0/QhpWvqRdP7DgCCJaS4OkQs+zGAEwbBEEQUyV54CowkRANw7/rFXPfxjHQPRgx4yYQORFGIg4pDEPxT7j6FuhpGMREMwdoCaalhACXFYgyDAM5CwlionwqHEpbIyv1RZJICIs4A5vzoQSFRktQLR3EFawykQ/xCCg5EcSBGTJw4KROAcAvHrP4Q7Eeh9ZAtmIFlQ3VLEexogbYYIRiD85AVlxMIPxiHPpnDA2s6oVDMhIU1CZCnLioy2PlQ9yBdecKaRmNUt5MgFdWgJAYPEgAcIQUKLFnJBjvjDIBjozlwNQgUofg0NptORMnKRXYHQoLsHmRa1LtSRLUK4VPsbUEgq5CCCePYjFhVIDP4x4gUgUyDYEMgjhHHhijSXp9Z8nWSz9gAVKEEXZVpviz2imDLu+MdXQitF2lKQBnvEGUBWyIAHbJEUDKGJML4eGtQwBTUYAxLXwENZNKCBA7TjH18uCJ2u9MlzblIistVIhyMiSwkrpP8V1ErzRRphDYE0QiryHMgEGMAFBvjZZSQVjAfCYZAQF3oBJMEvfkfsjBETBNGjMIhxpZKBDCwkCwLJQBZ0mYJOp4CnTRuBMVQRhwBYgAuyEIUGxmFWH2jgFZxo6wwM8Qz8EiS9SXaLkAeCrVw/KxJ3Rm1y/nHnBiWCpgzYc58H4IYiqPYFFggEHopBAYEgmjx9+IMitk2KgTjPGd34Bxj+YQRSfMIWe/kHoT9i6YocYSDb+EcWsnCEeWu60inIXjD4QAnOge6tRWvFDATeCj4IPBdYYMXhfM1ah1ZEzgKpWUqo1EX7IMkLy/CCF6Cal28dUCDaoojPCtJANjCjrUr/TAQvEtECXuzDEsxgxKQ5899/YCMc4/6EIpBcEGzcYxN/2AQ2bJ3ipcQb0wd59z+OwPSmiyELhbB3EGbQAkoAfASt6ARPO13pShciBbxIASVyYAEfL8TNnXlfVqYLW04pZyEki59GhCOQtm8kf/axgDLWxJxlQFUJnICGAgYfisH/IxQe6IHD/2GBWDxhSwrxZmCiAIJdBGIbq4j3EfiRga91ot0GQfS16YON/m1GHgIRw0BUn/Q2iMH1sOdHGwby7s5/zxLyyELXKz3vbfBjG3mW5w52QNKyl334AzHFBqCxAc+aHShsKK+M3iuS54dL2CMRY3et/w/SqABXAAhA/x044YJQmB8VCjA/NBDwAqgK4P3+aTwTLkD/C1BCBj04BCf8zH/LicMNECRfbnV77XZYQAFYErFXDmF6ZlRfENAGDxiBENgGbdB0R5A9X8MHhtAKAocGnUAJrUAnNWMJwJABYgABv/cPJMMG7cNaQVIy3MUZLygQI1cq1kIS/9InvlF+POgCHoADKBAJuyAOsRALrZALH0gJC7OElsCEC1N1lkAJlmAJBrBL/6B5BWGADKcRyCAQszcR9YUQJPAPJFBfyBCG//CFaTgQbYAMEFiGJIAMyMB08nCBGWAJ4sAM2vAPZSYSM4gQfbgUbzBd0xUSRmYyecYCgbALA7FQLf+2Mv8QcgLhAeMxHghwA5cACJrYCMXQCM8gDkOwDXI4EWO4ehahhb5WbRGhhgNRih4RhmhIELM3exBQi7W4CvyADNpQZlwgEL34D4zYEX/4IMF4ECIzEflTcYAoEDfwD81IAB3RaxYxXwJRIbtQeQghBxyhjRcBiQTRYM0YEW60EJ/EXR9wHq0RB3GQDQEwJG9gATbBBXNQQv/ggIyAEKzYhQKBdPZBBgshJYaWX+Hiiq5oEKVYixAohxBAAlWwC0ThiAZxWwORVRlBkVlhkQsBkVtIEObCKheRHhyRE/8QQLRlEIWIkd2xSiMiJIsnENxYjWeABWSAeauQB6sQh3P/eATb4ARkYAMUsAKZgAQVgARSUAFF+Q9I8A/9UCmD8A8rIBCDQA1X8A+oiI8C4YYekQcDoZURAQqg8A9fSQJ5QAJlmAd0cAXPEAgkRRDYB0rSGFNXUm2SmBASeUMd0RqciFqtZD8RoYqcsZcJUUqAiRA3EI4LYRsGUZIIoQO+QAOX4Au1sAsocAYvQJln8AHU4ApJ0AwDwXP0AAsGsZQD0ZRPmRFJQA8VgBDnUAFJUAMJMQiuQA2SIA6rMIcG0YUUSIEDEYG2WIa1SAfisIhjMJkvEAWoQwA4gAOhsAr/YJZ58ApcmQcKQALbUAhkQADPcAMMEm8G0YzSGBJw+RFz/6kRcBme9EFPItEAIqUQdjkRI5QQ5ICe/yCfIzGYFkGfGOFVBNEIwFYRYJQQYTAQFEANftkMNUBoqUkQ5+BXp7kCoPkPwgBcCMGZB8FzE2GhRSkMT4kBj4kCYRAGWBAGGIABhUkGN+ABoZAHzwkKNrmbcAgBjECWq8AICwmjYgkKV1AF6AmiAXpO1EAftbARDwYSSakDAEYQmgBGYtKeB7ETcCAN+jkmBqEKiABGRmoQ7zlPF4FQ/6CSB2ESByEE+PkQtEAL/wARnYEIiPBoAqGYQWqlNKAEgrACZvAPSSAMFYCAHJGgBmGhEQFcGFoQFbACNYCnGqoJB4EB1UYBjP/aqIy6BSdQppJKC7VQprVQCwuAAkY6ev/5D+QAEkZ6pf8wpEvhChjRXwlhqgkBEWj6D2aaEaowQqNHA5CZENBIEFLQqYhmFVYBoVUhqlLaUQgBB0KRChzyqgfBDY9ibQLRqQMRAchKEl61cP8QkAUBRlkqEJmAqAKBTJJTEdIwEHaJErqgC6kQB2PgBCJgquF2ECzWEe96EHrKpwYRr/UKWE9ZAcgkDEiwAuHQqwaRCQSxBQaRDapgsAVhaFkSrQphUwhBsP8gsBcRByEmBQOxACGGDtlwDQ5rEWbKsBkRaRHRsQnBIcYkEMbUsdkKYgLxAwJhB3BArSMRDcQargL/YbP/oJ+u5bItexDNsADOkJSpSa8I4aXfGhFw0D8ne7IKgRIRcbQG8R4N4Ck0IRDok65m4Dz/oAj/YAbh1q4E4ZoEkQQbYa8gIQxkixBJsALUUAOuUJoZYazgMBA25Vqu9RFJaRCQkAoWxbQIwbMFMbdQyxl5+7T/EAdzaxAUikEEgVT/wA3G5Lf55VcAyxMJ5VEhcSJO+w+sUCZwsF8CUXMEAbqp8Q/m+g8c8ghVWxGPo7q4EKUdIbkJxR4N0ADd4ATOEwK2YAtmQGhpGxFiS7ZrCwZQkBDJwA5w+1cDAVgaOghJsA5mGxErQKgCAVhJYAbJAAW9kA/58A+k8Ad0/9oPmlkDSfC2P7CsFyEU3MEK0oALOJsKd8sKPPAop2BrF+G4FFEm0gAHMNtVB7G6B+EPa9AiXnWunFsRgCsl/+W+QQHATEoQ/7W5HyEF1kqy6fkRb4drG1kqSOFxqKIo9SFeGzzC3mgQFsYRRqE4iDkUquITXiokLhISsCsQZPUWFXGMhfMPGtwdIDkQO/wUaZBFRDHDB5EAIvAP98M5AxFRQLFV9mkRu1YRlbsRi2cPpMtwOLyMgZgjpxGsKFQyrfosaGcQj1C7//DFBVEXp/ITT0CNUpEf1VAOKgAsIlODV8KAEJa3JzzCBbE+HBEXKTQRLREA7zcWKRGuPfEPFv/sTpgbES3pGw7zDxrXKxbxHAKSH64CIB+hKMMiA2PWi2PMx6IcEkQxOKG8EBF1IqmQVSB8EWhMEeG0xW4xnhKxlkeREDIrEGs8EMVWECWQCyFxDNVQXcVCEM2hHEaCEZisYQTRFTvgB+Q3yhdhToAszVlsMrksFS2BvwpByxuhjE3qEcVIEL6iJ7CiDDPAB8FACbFAL5Y8EEXiEW9XEAFQDPUsEDIRCbUQCaxaEE9hzwTAIItAAdJQzR4hBekxAWHVgtLc0AhhDdksEaLyII1MHolcEBBHEOpJC6U0KAPBMQJBLHvHAlK4FOXAJAlRzrziKhFhAURwA6nQyD2AUeT/4RAVfTIezBmlVSn2exFEkVkCtMPUIpHPEq6p8AxKLBHlkDW5YCMsPRHKMCRxvNRO89R1EtLlEAiz1glUEAjPoTF8EV3z8iYR8Qa1sJ4KUQJ51hHc9yxS4gMLsRN2cAbE8SB7uBFuTBGvzBVFMRA3nRDqkBAOO8M+8Q2DSx+GQxCk8Xj/sCWEQAhYcFsYgAhC8AwqUGVIgxA4ogwq8FYE4dEgHTEaCCxUnTCG8DoG0EcDYTBbUzpvMAUj0Algo0hPFgwzINsI9i+GQDWQZDEfrRAA0NYEgRI+wwcOfdzIPbHE1pbPMgu8QB2CITfHEdLBAixbZRCEMgKebSchJBBV/wBX/AI8y1MIVIM8VbADRJMQryM7AkE1wxPezFM7BjECfYPas0Ldu0Es7VxJgTAGa7ASRFwRe/wTNOXHvsYKdTYQay0SrTw5EY0QRywRf004vwhBJfA2oWNtSmAM7mLcB5E1sy0Q3bYQ3SsQvcAO7KAIZqNYw0MGtPMPt/A8BBFD/3CP3ituBHGPjMAOAiFzMbA2iZQ80TUQ2m0JT2RNQRALABIIYiLUBkGqBqF2BmF3BPFl1IcRBt4RXwbXGWECeAciFiEUN2hGe90RGcYpT8wpbMAG2sAM28Bpn+Zp1jYKuhNN2IRNHi4QVNYDn0oQiRsRm8tCuFBUrPA3HKEIIf9QQ2NwC2OgCCTAWIwUCNazSNnTWJlmCZMlEIHQqgEwNJNTXqVCJaM8jLn2wEg8EOMsEUzQAxzlEaCCUb/4D734JFhQg6rdSLje3pLQBIrwZENQX0MQNnwDLH1uESvUuAXRPwyIxxNBBlcgCc8V7RmQPGzTSNdEMRaDGqpFC8VgduH0DyiZ3OIeGvppxuO+EUrgaF7R089C3tR+Ebf0VkvNQSWQA1ZgBeE0TqP8HTpRKU3xyAXhBFfSEw9+EQOOOGsQpBXxYNTBBzx15wTBT/xEESz0Y0oFMQJFUFow5ueeFYf9Eceg0gJhUhUBKub08WZxEJfCBO6S2AdR1xFhUlH/3BH3U8MuJUAivBlqVwVgFAh3wAvYRAm2TYUHYVfiQDKJZUvi4FghIRQowc30YU2LpE1x7AUqAALZELP/YA8IQVPO+g90Rx9hn0A0Ea6tAQi9/A9L4Bk23/E/8w8ZTRBZ9iCtbgyUwAIX/g+twGT/MFezmZTvsLjERRAPShLEVQPNKE1MvxkT8zbNAQAk5QctMBBc8GEaMeHrgQMWiypc7hFpvhnPd15AAcybYSUHLxW2vBkQuUFGYxCfJkSSILH/UPjnTk1ocNqTpXHl0HhEnRBh5vbA/RM2j9YZkRbTZQFBMoxWAuoJkedSkfMc0cP/cM1beLedMXrPwlNUYAAx/+Y25WAaKkAINlXwk7MpG5H6iGP+wD8R4BWsJvMD6o4Q1voPV3xhfG8QoFdEn8ZT3A8QQahY4qOmXLlASuCowvMPwT+IESVOpFjR4kWMF+f0mJLR40eQISECEPkPiMmSKf+1+LdI5UuYMUsCkunRDcQLMiZOYPCPA0UVIWNAdAbxR02LR5EuLZnlX4YMEDOkmJrCgFUDBiyNmDIlFo04Al78EyVKg4Z/Pv61gyiLSy5LXIR88wgpAlO8efX+c7DXb8QLfwWDbDR4IgufPLkwWNzCjYVAKl5ArmXDDMRNKTEYFfypoue/USWK/pglg2moVVOkCDJjRpVf4AQE4pIO2v+qf7z4xJrBZ0ar3jOCPRt675+qf7oML78YxeObfyQb6pXA3Pr1mpEiPojo5V/hf6g87viI+N9ixYzdYHrzxgIICzsCsciF+x8S7BPtbVIU0VaMd/55BBtswgEjIkU+6QYbXPByapuKnKKokH+O+CeLLI7IQp4stsHwtBQMMcSSGUZQYwQrTCyxxGCCoWobXgxphQtj/nkDhPxyVOkL6HSMiZN/gGQjyIgsuKiAw3yEaAfy9JrkmEkAkFKAAJQILxQFJpoDoycyMgUiniYQh4tVuGBGHqj2WW01SnDL7KK7itoLG4hwodMfiB7Bc6IGdZQHIgvFkOgIMY6wsI1/Cr3/MItcgqFkn3/2gYoqSqEybQguWPpnBBwhMvLTHWKhaJENrhPyHxf0KlXJmmiaKCiZKPknFyVJEkyFHEx64AEAAjiDExdCwVIBBbAMhZMXqBRAAAAEcI+PJ3K5QNpKnmDBD04YYAABbRmYwA8V3gDgjR144SUXPoADJoM/JXrTorvuYvUveQSFyN6IkJEIX4jaaAMZf/8VONF/5LFExlb4MIQXeVZJZ45XgrzgCSae4GoHFeTbYYRYLDE3l0PEgQbIf4acqMfBOCF5ubH+6fQfneYdrEtWbbVOi5MCqIMTD4QNBRWfPUAgCkJiqSKXXGLpQYVY+ED3CadZ6KGAbbjQ/+bqWXihhJJWOmkF4UejyoBCCSWy4aN4/xlqqQAHEwK/fxih0C8I/oHgbrwDboNQQzPMUB4LK+TnH2SQgaANCPjZRpxZDHGDC4mAXFlmyiu3XKIuZDISrx4kgpUiFzwI3YNFbsCjkUaK2UWcXNYlFKK67a4bN9rtRrSiwCMq2y8nYopgAYrkZe7222Nfqu7bK4zIQn0Rxfv5VbIwk2TIkcryo+oh6im/lv/h468tLIchIpQ98oP7kHDcJSQcKgIEkGvieL8YZo1ZpfB/7DMeAkb8GuPyiQAPgCkhQUUOd0AIrIIEhXjGP8TBqvXZ6CURLAkKIGJBmQXgHxrU4FIuQf8RY0ShRv9wzmBuwJwvUMQTEelcTEiSwh0UwQLNQgEhxOEBh9EBFPaxiL4mJJF2/QNCV0jGLQYIkSRghjkFZAooIEICKJIAb6Cowi608w9fCGA6liMCRdQRkQTgBYNH/AuOAlESCsjkA2kkhCdo8I8rusoiY5xXBzsIR4jUwSO+8MU/1hcIECgBBWHAABKaERFnyKkZFfiHMP4xCIr8rySwsEgNZOKKfiyPcPvapL4AlryI5AEUhYgKKHZoN1RWJA8UceJEWvkPUdKBDvGgZQJCgYMqQEQFUeieRK5IOQJMJBT/GCZFsAARPr7kErugoEVK6MdmzisOFCnGRORYkzT/SoQcEFHCGc6wHGsA8JcSCYNErISINyLzgi77ByEgcgMcuOIfRamAJWGxAno4khr/kCdEIGmRFUCkBjWghx7+cQ6lxEQP9IjICqjhCiXQYBc6wAIGcHCFPKyidga8mxQ9CoGP0mEVkgjEGRKCAhTgwRffJAQGjunOiPQxIh+MSCb/cseP2NQi1SzJPj/yQQ3WQiaBJKNfTvARQeCFpxEBRDgh4tSXFEOmEqEjU6bJDeFZ5Bf/oAUW/6EDFAgBIuWECAUogANqrMCR/5CCTA4Jkrd+RE5JrEEFVrAFRPyjDoIgRx3CEAaz3oACNyCsK24QjhuEgQa1qEUAfCFVPlZz/xdKoOwZ/4GC9V2CBlbS41gh8s2XVPUlfexjV1NCC56aliJ1CN+8jvqSzYAkExNRji7gQJEGTGQNEYlGRnY7kTRcAzl22epfAgoRg1okG4DIxlKai5xs/KK4E3GHXlIxTYzEIRXZoAUiTnCCLcQzCZZM4j/WIRhGLkUYKzjuOoSRCVeI9R9JhchsY1uRE6iCFtwtBi38q19aHFXAR92qaj3SXANb5ATp/AeDM4IfAZYkoMctiSYmQmGQIOcfzYWIhq1UEQ1HRBWqQEeIBQyRvHokFf+ABIsjklXgSSGuEbktbpeS239MYyIr/gc3ImKHiPzgtRUpbiqyep+MQAIdE//BrkSUAxEdR4QVFYFEiP+xZI/ATSIR8PFHdlvjf6RBIrdNAyvgAIdNsKM/ELnMRGZbXrykdyKMlPN5KcJIgzLSzkmksDDOK4waDMKnFJFvI3d85YqsOMSqiEAq1rYX4d3luhGRX0UikGKI8Fglml4OTTh9ER+DIzmjxm4EWtzVFvsotzgWjJgj8g04POIfCeVBKhJap3+cItUQEd6t/+GPKfv4yRGRRkh+G41iT1lHDVjDqr/RgAZgwwxr/oMtLNPm2VrkzeFgRC/+QYp/JMMG3fgHnCVi7vO+KwlJsDNTkrgJW7ADIr1IhghcUQNhuGIFM5bJilMxZU5nlQeC4TT/K2rNiikXOw7cwO6nL9In2k5k1yE5ZCp4PGmJNJkiLYYED3xc7H/gIhrKVo6yPyIFOTOH1Ui5ZlFdXhPxvFzmM6d5zfMyTopMQiK/tcgyXiJriHQQEF3+yxbxwuoU4gQi44tJMf8Ch6VSpB5IWYJMohwRHVSdIsf4hwAscsx5bU8vHRCMyZVk5YhMIO0y2S3PU8J1kZxEJdeASPfuMBivcwcmnYXIqm3ul+pERAso+QfTB5OrvfRlgKP4e0oQ08KKqL0lDxEJTmGy8p3XxOsZSTpMmA556+wW89chwiFEgvhcNSkQkGHnLqoJh2b/QxJhhAjtt9R43OceLxqPPEiq/4EXy7/dViukSCRAPhGSyP0fxCdjbzNCM7KT3TDSh8gzQeIFTOQcIuWYhBcmcZApMI0IkNvF73VvHcqfPz8wCHzwS/IAL1TDO2H+R9vr/w/nX6cIEQm8ReoBZpm4iaXzEbfLD51jFS8ohxGQgVawiJjJC63DiAYZAPWrQL9wiZrYLbr4B2/wiKmLA5wDj5TIBQIIpomgKb9rOcOYKsvZvItQAGhgg0PoHPM7QPP7iHJIiQNUCQWkmX/wwbwoAYnAg4YAOgvUi/RjCg17GZuzPyCzmYtoAN77jpRQvi6aiOnwO+xYAzzYv7wYvZKAwongBFHhQe9gFgAoh/mziBuECP9lWArvmATyoJWIwMBU+QcPOMKXS0Kny4s90Is7mhyMKMCJ8DHMG7brILsk1EPmkIN/8DnNA4AdzDllSMBJeEO9yMGR+Ice4IKRiYg8hAhCXIrsabzYS4n8Y8SIWJWU8Dmc+wjk0EIRdL+8+D+ISDCIMA5WG8Wa+ByJQIBiup6XuEKLwDKKKIGOWApNPIZq4LplUMN/gDtMxItl0Dvtc5lDUBlBZMRFNEGRiKYjCrEXMDzriDm9oDuI6DItjAivc0EwRIoaEyobe0fmEEbDeIPv8YhKfMNyeIAR6A01qAZNtAiSqAaSkBIAyD6JmMaJgLscHMiG/Afv8AJleEaui8P/G5SSf3CDh+AEDEwJJigqsZM8kQA9vbhDpFiD6coLJIGIDiyJqWMKF1RF69jFv9BESPyHHFSBRrEEndRJ7+AO74DIkBBKZdA7TVzDiTBIhGzHXQgAKvGFACiGXwIEXYgDrPQFIiAZs9OLn6g5FmDCf+A3miyJPlSJApyGD+NEm6NHyvE7zDOPj7AAFrAsHPTHWKACWVFK68jJiIBGi4BIwGRHTxgAAjgFkAjJssyPs1xMi+DFj2gAV4sIWsSID/AyC4TLlFiDbLDLimBIiSiHjjGE7UgJvny/f1CGcpgCTXzIiUhGkOgBApg4ijAOEpoXI/wIsaucYWrM61CLeQHA/5oIAOy6OpmjviNyNSUwBl/0iNXsCD4YAaIECV7ZPNeUCO5wTX6EiAdYzVgIhn+wLH7Uu/BjzX94ANjMCFx0zJRATI/AsWgALfbECNsUiYF7ieBzSwCCKcGwB6AICR0whvT8SYtAz9UcAUM4o+lcyIq4zhwcAe/ZvteEze5E0H+oAkuwhAHljhHoBBHhin8wzwWNjujwBUS8v4oQQrwAAWKsQF3whMssifpkCuREn6XYwJDQz49ozM1pPDBUUfyCCFaIgGewPogYPOVjUPT8hxmIiAFdyOwcgWAYgfmbAjUATxHR0IFczWAwBGPYgYOQUojIpSAIkU1xUgglTQMAhv9NWVDueNOReANf+C37y8WIKAEglQkaSLoW1YvdpBzfHKC1pDkcnVHsgIM4iLqKOJ95uYAOmIAW+JZv+Qc/IAIacAeuSMYnhYiTsMYH6I2KeNMpEFUpNYRg2IEpsFA0QIMqAIYhyIURyM4paNJ/SFBfWB8RgQg0AAZgkARgyCUqQAMmHVNgSIEmuNBgUINRPU9m9VSdrIYdOANaAAd0+IXo8oWEuIvJnE/DuL2KYDUd5daU0EUfMVSMYFQlWYISoIRcUAEIfU3U7FQWaFLueENHYE0prQIBVdUL/YdgpYIqyIIhuNAqCISusNB/EFZhjQg0oAIDGNhbkIQhyKWJcNj/iWDTTLVSuHhXN9y+E9E5kpiCM3qGX9itbW08IHu5dZSISljMcLW5OFAFEXQ5yYPVf1CDf8gVX1SD6IQInJ0CINDUv2Sad+2KKaiCW0jaKuhS0mRVYR0CSWiCP/gHMACDYB0Bfp2IXR2CIUjaf0haqKUCKoAIgJW9Y5WIJvDVUqWCdRHW9MxUBKXVZwiEYAgE5Zg6OKCpl/vT8xNAH2kSAGrDiliDOBBLvciGBpi6l3U5LuACXjCRigAGBKBYiGhAijhYiDjWs42IKygEMJAESZiIEPiHEEjatPVXXa2CKnjYIfiDJjAi0u2DWzhWNqUCrlWEJrAFieiDEOiGBcCG/xioAkmoArGdirEFz45I1U74h2DIBVM9mirwBbrIrZjMCNGCCbZgi8tBiwM4AJXoggQwgYxYXIhQjs6LCDo8InmcCEcEiSVTyOxijnogX5lrAT9AmndVg1iQhAWIARSIBZydgSCwiFTNhdediGS4glCKiP4R3dgAhwXog27oA4mY4FH4Hx6wAx6Igd5ZYIloYLOJ2HUphIGtVfD8hx0whk4YWwNAA0PIxxEwhj74hQapXoy4hJOViK+cCMOFCLbwXrSICQ7oCbB7iSDGB4jw3pfIHIygXzhyQaYLjL2IGCauCWirRXHdi1loXEtwXqQRW0sIAjb9BzKACHdQXQgdW//mnVA3MNGSyC1c0AWEiwFw4AFdqC2JsIM4VonzGoMxIIMhyN1/GFixDYZUBU+HzQADINt/CAIDiIU32IWt2sBIOIlNBQkgSQW0y+JS+IcuMAHa+9YsRgq/tOEBgt+XWN+9KMUBECEIxVo+0AoIkd0maIIhGGN/NQSstdIQZYEGUhuQALoTzYsMnjIeuE8nKITQ1VU0EAgDABFFHmA1DtEL0gVms7mP9JETQkuRKIzKZBUYKIEHHOWJiISZhQkWHIwJ8IQRgohg0IqJsAVbSNshMAAqSAF+OALK3ZRggN3LIbcY6K0mUOZlDgKBoIpFhogBRt1GNuSDqIYoqAU4qIX/HXCEmfsSJXEBlDQ2FJ25KibndrKxKawIC+jR2HQwmLiDcb6IOiAHUcHZfJQIYAgC0EWGK+hcZEgBiDDdKiDNE44BZ3g0jAAyomaFlKUIOZGJbiADRQhdi82AMU5oiTBoieCK7oQMAQiKwQNprr4IUaAcrRtQJ94LMdzbilgAQmhnkDCAhf7aURsDobYc5fiFIciAgYVqqRYJNOiKBzUGNbCCfwDsl0jFLUQKtVirL+zorrbisV5si2AAQRA1kMZllRjbTjDkUZ2CEhgBLcgBLVAD0PQyiPOLHdatmNDef2ifvcit36LN60jSmRPOwShFmeM5lPYIC5LLReYFpjjq/yMUiCC47K5ATxYoATVQA9h2bB25opl0IUzwy+auiEW0CC9kijKYR8gMia/+i9C2juvVYRCilVjO5X9YZEvIa4ig7H+gbPVGCl24T8uhguB2aO8YgSUAgl5RbsqJbsNAC1FQbbdsEqPL0chU7IigGb+liCr+aKTYvCKobt+6BI41DJcwmX9gBomIUZ90jfO+2IjAZTZt672w4wweIPkW7n70AhUIBOLMbv2+DsSLCZ3zS4vYbonAtOUAQpl7ARnqcZOuCRvfi56mAl3u0ITW6axIcmCgAB2QAmdYgAj4gR9oK2HYDFcwAzJQbcFAb8MQ8YgwBCrgCi8AAIimBTvIrf8P44JZgIjSPqI//IcyzJE6jYgaPSILUmWJyNPG4zsXMomx6J7zlYhw2up56YFcSIRN4ZgyzetFXlNJ2IQG0RPssKQagIVACwccIAOdVhJpboURMD8joQUl8AOS1B6Xk2IWCPSlUOJBfAn+HoxOzggpVu4Yp4jkdrlA8EmI6A1dj4iBdXQpeIcfSK6UGF2YIHaGcgUyaG8dEVs0MGSDnIQioIQWaIEBIMn2lW3B0PIXz4tYr4g3N4xZXw5B7EpVXMuxgLwmJc2JuApxkARhIHYdYagBamsXHoEd+D4vGAE34M8c4QRuP8Ky/uaIsMfB2IM/DIxeqohsVokfNwwG8Pf/kBBAcgQJQvcR56iCmPb1ZS6EK2AEdsiks8GOTZAXC6ucTZcIZzeEErHEciiANccI1F4KVlyONbivkAhi7DDHi+A6rlN1lZj1ZwJciDCFL8Foj0j4ytHP/SPGBI8JtABOw7BLWimEbVjmj/A1XBsM+GaVEp4IgQjWVZVONZyCaEk1Wuhh3eOEUoGG5RjwblcSRY2JVcthpsjTSij1mjiKI3MXihhtcS3hrBCIZm5YTz+IcugBGliDNaCF73bszcFEdC0qb52IWdfzuB9AO617iKDxmhCV61a6mGeKtDGKuAa63PSL1Ef5f8AKR3b2TpBOL5iCHlgboFfuH9cUMtro/8xnjoh5idBHir7v/bV2fWCQb11eTRV4hicbiyCe+QFCi+bsar3Pi208ortDCtNbYgZXCT6oc5lYm+FPifGfiK6fuU1XjXpma7aO/a4wBrD4BwvggrM4i7W4f4jggkR4AnIAiAjf/hEs+M/emoKEDDJs6PAhwx0QJ1KsaLGilosNgWjsCNHUBo8iR5Is+Q+QxzwmCxJhMIEDAwYEBywcGcPggpUGb+rs2TMDQaBDMqQYkiKFgaQGZqiZYuzEPwEguIgSpUEDwXbtCHZhsK8Vnyh2fJIta5YkDoNAipgccfYtXJ/ZDE4y+6SgjH+H/k1gwMUvgwFuLPyz8MJCIApONv8hiVvRRsNPpDwaKZsiqMcs/7Jk4JyBaFEDKQyNYBELXBypOGTJqgol3RxOiUrwqT2Dz7ObDRrY+3fPMXCzAswWeRH8uEl4yB1GMuilIUqduQqW+OcScF/BxQ0jLrbACeTlED89/JTv3yfJ5CcXJO8TKEHNGuVzrv85BWhLwfhQMWbMrVsqjDDCDDOUMEMrCN42gyGE3KQLQW+IN6FGEq5UykMSULghhxdF0twk1RT03FksWNfXXxMgINgXFuxgAQgwgtADJwUJ0eEjDfjzB3mfKLLAI+88soAi7hnBzh/O/PPOO2cVYpE8BmVRSBbyTJmFZ58ZYEgrlrhFkBpMjbD/RIF8IGhICpTUZokxtETXIZxxmmQBAHiQFUhB08GVgJwELUOQF14cI0BzCDhkQkMiUsRCIgVx8eg/XPiRSywquHhpD7FYQgIFBOUUHDYGPfKPHbYY1I1B2DyCTQg+kvdHDP74888pJsFH0ZMEHcHQrkdk4SuVWAqbAhV88GImgVaIOYIhVBy1Twby8JILL7wUdm1FLhBkirXH1TghCBIRZGefDwFgkLgm8fFPdXB14ZGFbz0QqBfLEIoCAqHoa1G6EMFUEIqraMOFJYb8UxsfsfDRSi7b/DPGpwRFABwuBGFT8T/YfBOqP6M2uSouqjLUJHBRRrlrQ7uKccTKLbNc/2UWBgRjCC/78HIUaEfh19lnluxDiYkQ7RBLC3Fywga4IERYLkkceLSuQU/00BOGJbEl7zLLCEqoEpxAo68CChA0h0O7nGuRH9YS4UcHuQQizjbbDOGwPBkwI48lfGSgUkM5TdzhrP9U/HHGhTummTxiFKQ4QYz/0wbLR0DOOMpHDEHFDFRE+9lQn3mexRA2/9OKQYSZvkMgO9zhxz+LcMKJttZNaIoLphAkSkFbMd1hAGRV8k8Bcp6tKNRlTfGAMvUCEMkZnOiLStgKhBI2J1EMJ4AA52JiwbrB//47DP8w81dME3AxAC+WfgHA29vwM20rNDsMkRT/1E/hqA+FCv+c444ThMwRkGEQMbSBgAZsAz8EWMB/pKATM5uBJTZXt0KE4hWv4MQTLqBBCVzqRTv4YOpiwYVt8IILSCMIA/ayHKeRpF+7K4s1vOGT4O0hTmd7yy4YAoRlPAAAAWje86QXClToCwEvCEAABJDE7O2ADxm8QC6gKANGxaSK2ZGDCgCwg2oZQkFosESULKIkiZEkfyIx44QEyCuKtAECbXijG93YBmQAEIB4M0Qw0MAHNHSCF7NYhfgoQYlc5IIFpuFDH3mRAV68zxC52AfSZnHCCTQkXHGRCQtbaJEeYOIhPQjfCz3ihlBSKIcECZAylPGPANTBAy4Yor5g6YIBHEL/HCN4gwB2kb0ixEIGT3hCAYBZgh4cAgF/QYBf2BC3aS1sYQxKwTY6849cGWQMYvzH33risSU5ZhNkaYND4tjGccJxjpFb2TaOYglLUMESlFinAXhxN37wA4FtkAcw5PmPb+2TIFwgJVmUBtCB9oQADxkOXHKQg39MgSCe8IAHQhFRfb3SAzgAAQpykbDa5IISLajZLPaxD22IVKQlTAQvBCnITnSiFVRQJHzkY5HGEHQ5aoQIOCcCgYK8cY5iUCPK/oGyApKABKA4agL5IQ5LjHAVnNDGNubAhvM1JF4d2cENa6pVu3DIEwhFzpe+8A9P/MMF5nClC9LqAg/IAQ8B/4jELnLBJV7Igx/b2Ad+eGEAS8STF5bwa7WgxQx+CNVX8bkVcv6w1X/c1CDgzGlDIKsREuwUAnLUlVAVBzkEEqSylrXsOG3GjG0YylBksepiR0KEf6w2tQ5BgUAbMgCC6Mm1BqmJQTywCA9wggCXAARwG7GLKogDGEcIYGct0tigQiSM5YrYArJJxp7wzTEkMAkcP2vZVUAAGdtYxTb+yReC4NYgsbXIHUiJ2oJE4R+jrMgrNJKWhtzAJDL8hylJAkqR1JageCqIhi7yW+ACwhqNaEQguJCBXQFyp/9w8IMp4j/bTuR+yIFwSa5bEWTMcY6P0+4q+MEFccDFAwVBwf9i06sRPmmEAgbFAJza65D1AnS2D7HTV0uCEkDEgcfZEMD63hCLVRDZIwVs7ENkKieedKQCFH7IOLvb3TYqwBjZi8pD8mtbGjvkvMhpbVzI5Yt/jNkgKH6yRd5ALtSmd2oTmW/vCoKOf8z5HwDAxPYsYAEBBGIIdKBDHgBJEA1TJIxRopKuKiefcDwsYsgJT0es6RMMW7cgEKBsd5EBAVCIA5erxHJw7CRqLpeyIDRAM0UuURA7qfofz1gJAfDUA2OQRcsFecGpyUURW4+1ILQWyZsIgj2CmBIFH/jHDQggDnF4AJB5oAMgNS1ADhfkCIV40rULsQ0n/MMJODCDDf7/EAIn9CMJLxwEowkiggczAiJXICUoilrUSxe1CjvAXnMK0mrg7ELUqP53JTtU3oIU2CcCGLMuy1LnguT4EmStiC8C4Is3PMMYVSDEDbbg5HMUZOPN+McYa4AT4Ihc5AQxOUQG0Y8rUNMikiXIUf/x7oYI2iCEfkgebl6Qo4IiDz0HxSvygIBXq+C/Bsk3RRaiaziZo6v/CIRYK/IBAhzbIxBaeFziDJF9T2TgcUHxqTuyC61fxMYVIXtBIlGLM/yDEANXAkFooGpV7+IMIHgBCM5AAFc42X4gJ4gzzqGHf6zAJLCYyOEdQg96FD7xEzGDCHIVVMip8Y2Pe2wcLftg/2TQoRBj2AU5qpAvn9Oh5wRZRbsJohJQwLzdPn890Okgii68QgHrPgvbGdK7pfekU0zLPUkIAWOvO0QJcTDL8Q3SO7T7xDj/MOiTbzDflegA+G3HwtNP4Asa1MIX3a87Cs4Q/irgwBXUWEEFPh54Yayg8AUZBEHgrxHHwyIJSahA+gnC8X983CHn+PjgOYQruMIW0MAuYIACrAKS8RRDfBZlPSAEXMEVvMI2YEH1ncEZvIDdjZ0vKMHFUQAhUMDUVQH2/cMl9E6ZUUQd/IPzmQTz/YOdWJ9OQJ941MI/2KBZbEFBrKBZNEBZwJ1IkMM/nFlc2GAxMA3SEUQjXAQiIP/CP5waDt4Wst2A+dED/+GfHkgB+/1DJjgZPdRA+/2D/BXE4dUAPZxD3xXEOfzA/vWEMNDDAAoCDfgCCmCB8IUBBlBAs/kcI7zbu0kWBAbivD3bKogDOewCIhIEFmDfQpTgQ8CYR0RhRxSDLxxhcBCfSEhiR0AFwHVE2OmAqR0HOShB2DHEfUWCNciZRngfQ6AAEJKFNRRcQcQBJz4ELdwgQfgC1xGEQd0ABVBhDQhDOAyCMIgEx1nY31WEM/TfMgLeP7ThOYwRyCEBGNIDBQhBLdAAOQhCGHRjGFCAOJCB9I2jDZABAtxAODrBFRAZ7AUdoAHa6xGZB2wDBtRBGGD/nyM6RClaBArsYyYSRDFoYkW0WjH8AkXAmAyShEGKxC/cokeYAUG4wj/cyFbVIlTUIpykYiwSxDX8Y0CSWVwkH0N0JEcahCoQhBN6yhD+gxKQAwWsQDiYATVkQgBu3ESkoRqORP/xX0Hs5E4axDm03xnWAAZAhRIIgiAQhCDkoS9SAAW4wlM6ZRhwHy3UglVeZfdlIwpQ5D+AIkFcAkXy4D+IJYfQQDFYoknMxT9UpVY5WlwkJUGIpEbAAUOsAV1WBDqcpEOcZCqIR7D5BC0UpENOiF5SRC2cAA0k5ihQoUHg5EM4pkdwHMcpyWQWhDRSRAUkQTgIwzpUAPtBIkEo/4EmvCKMleY/wNgWnIA10AJrZkNVsiZrIuZF/gNGMoQmQMQtuoNG+KOc1GZPqKVJIIJeemVB+Cb9OMRtFkRynkVCNERCrEFzQggk/ENKQsIt9qVB8EBBuOUJqMJCPoQO/sNyPgRwNoRI3uVFzEV5WgRcikQapME/pAE3EAR2MkQcqEIqqII1rAB4mFtqpWFn1sAg3N8/rMMmCIMrZIIOcKUOjOdDoEM2rOc/6KVBGqQTNqSETkRh6sQ1kGRxquRcbGhJDGZFgKZDGGdDiOhKnACJWgQkYCQydsQ0/IMPdkRzMgR6Qsh0/QMrFESPVsR0RkCLmsVY0CV6loSK6sRYvP/nfEqDQUAIHOgCHGhnuykCQfgnQxTjOvwDZHZEMRLEl3JpQRQjmf5DmFaEMNSAK2DpOnDmCkDkQ2hCJnAhnXpESk5Mkn5KjDLEnJoEdk4MoGITfcYBOsRBX9anRwBnhmqENznEfJakSFxdX0YAIgTqd1aEdmpVNKSBHcBnj8olRUxnQWRqxzHEp0RAoNIZdiLqRfyoRwRpY5LEkRbENCQEHEQDQUAnD9iAEyiWYnEbyqEKyjnGmZLEOoThmBIEPSTBCkik75GEhxrEofJEncWAiKrChv7lPwSgmZqkqHqnQ2AdRPQlOkQrSUxqbaIoQyDBAogqRTzqRLAqj6ZCKjD/2S8kKUHciDchAU1VRK0YBHxCJ0TUaFk0gK3CwY9KAy7gKn3Sirs+BA/8wGUyxA+kwg88hEjawVjoKEMMBEEwLHwShJNaxMU6RP9BgqFSxBr4oMESRMv+A3Su7Aqwwz/8ga86QbpVRDfYQDIkwz+EgDdhqUEUa5YWqNB6KUNsabdeaaP2AmQMQiYMwgpgjEcc3/GBg7T2aI+y6sVqZwzgKUR0qUH8K0NwLETogtkex8M2RP3IK0mwAl2G7D84aY/ygHZqp7zuqUVQrUawLI3GBcMaBBw8Ai7wACsYrkPIrUUEjuDQWUHoaBqMylhYRAPMaEmUrE8kxDc0wHfYQAgQ/4Qt8Kr7VUTJdYMTMEI+9AJB5EPq/UM4rEA3bEKjFq25pam5Ka1GpCmqXGlBbEI4MAIU/EMvTEYyiEA/rEASqCkFrG2kEgQrQEiPPup0XuysRIB2gmrzWgQrHK7Ipq1BMO9DcEN99mXJuq1HpIKhKu5EXGwqcIOOzqjlji3AxRkgEKydnUtWdaL+/oMCoML+/i8ABzBwJGFD1IUAHzACJ7ACo5m2VsQSMsTZGDBJNLD+8lNHqIBJiI1WmRYGwwlHLDCF/Q71AYfAHscXtCBBRN0DX8TIChtBDClZzCpEhCcIk0WO/UNGLIMa/EOAjcSNGkT8OsQN+4QD/AOi+F0NG/8E33aIDGduSfxwRxTBDh1D/lZEjUZdQajYWzSxSdjvPyzqYt2XSNTXQ3wwcnQwAAwxSThAERfxC/0GCJPVHaCwbE2I4lIwRQBBB49ER1YxcPwJSVjw3wawGlsEJqjAQhWEHhdE0NiWGxfxESdxKPVwWeDxRTSASErwIPuEDAPAMRCEFnvEEvCwRjyAJG8yQ+zwP8glEp3EkT5rQZDNKb/LSJhWuVzNKUNEAKxwR8zqC3rEL2OsQ4TyRVDyWcTOWaQBAQfHHVRHdQRNIIxAD4xAFBgdim0fCsDNKmgw//6DieWySMgEOC8HJfUJAPixThTyuXwyKFOnnMROKDAEWaL/skgEs0h0QJ4QREL+A4n8gyb/QycBSkFUwySkkgWogBsQARcwQzy3F6mNM3LA8kSgZQLbmC1PRD8PLIV8gZtVBBePBCh1dCjdBXAEz5fYWUHckKKsxCR4wRRMQQ/ENEEk8nKMckHgMkNEg4lCtAKb3UX0cxN7cXDckAQY8/9CMUXgc/D4hDhHRIc8RzkAAQvwQbtYwXGUQbtUhE/ztAJf9EQswyT8SSR8NIWEDzE7BFmDtL6RRTxfhECyhE6IDTToxYjUBSDHBYm09D8XRDlMwhSwwAWUwEnDSQOgkQA3tWvNNZyUQ08I9T/wMln4LUGkYgqzM1wELkXQ4Ergs0Zk/0RF8AILqJJGiMgn3zVGjwRjj8g/PMAIBM90kHTrFMQijISWZbVBUDRXdwhsL4dXe4RjkwRk5zZwBPRDKDZBiMhzJDdErLRIPIdpe0Q/70BeFIShnJBJNLJwZ7dJyHBCoLN99s6wPbZ2w0koMMBZH7dAQ8RzWDZF7LVPKEPQzIJDhIRP8N54668YG4S2ILNIJMRv37dBiPZEcLNrsTMSBcA6P4QmI7dq+8QOhI8gk4SJ2DSAx4mXLYft+IT6gvB0s3Wc8BBqF0Qx9E5dZLRB9DVBpHZZkMi5qAARWLdzVnhB/LdGP0Rvl8W6XMBbkN1sU0QQOwRShywWI8eNA8co7f/XRZjxQzQdgQMHTTO3SWjPck8CYxO0Tqh4QRjw2QBALnAAGywCf8PsSJSBAlvDjdYDSeB0j5+F0hAGQP0J8kwEvNb4P1D2SmQEYpOFPZuF9BREW4+ECtG1KfYEiv8Dlqd3igOKihf6oTuEezNEPwOyiZ9LD3AB7JAEhdN5nDBAJukEjT8ETseF+WqVDM+nqu25eE8I9mr6ccQzk5cEmFkEbaiyF5gyRXgBYzO2Fzx6QbAzJkxCJz3Hrzf6P5R2iJT4n5RDvTAEnK82RUSBOHzLbnkEmXd4RZSzSNDySFBSnsv4CyF1Q7BsGth5IZsFHABCcD9EA9igkjvGn/tEoEP/xBNMAWOrErGf+ANMQWncO0qDWr8DQLITBK8bOpVbRKH7Mz9DcGH4Qbd3hLU7RiSbRMPDyZr3BBGexXtNyJAD1DIzxKcbxMMfnUc0uUks9UQ0FEEIuEHYOkGwNoLEwhTgeoMbsKKQCEGvdJW7d11I8M5bBP6mtEEMxwuIw5q76kWE/D/gNkFg+4Q0dZFDxB6XxQBUvFaZfEFs9e5Y8nKAuwKrkjI8t7OXQzmMAB8YQrOoAXNndF+LCL+fOF8XBMsfFBJFwi4fGIE1QjYAgrgWRILJxAe0sFkwvW1dwoavRJjXlNUTxPTFM8kbhH07htYDVOLHSaOUckesy3SYuKG//32iv8VzGDAmHAMm4O/oV8PZKFGcfUgAYIF4udbHOwRxVsQTdDDgQ/Tj+/lEeLd7TgSq/1vcl4Wbd0RWMbYZ1/vmF8QUzIx6N3jCw0Vy57qzn3hqi4gyTMIkfNUHRHhZ9AWqFb52D5FJcD3lOsSqB0fHb1X5N8RdAoIAqAALpDa/C/gDqIEjGYJE/D5ZmHKj9zPLA8SyBwK9/PtXzuDBhAsZ7pDz7xRDiQZ7TLSYcMJFjRs5dvT4EWRIkSNJhiK5ENCakw1OJqzjqeXCOCMLxFxpMA1DIhPPJAQEIpaKiUASIjSo7OAIS7lGSFxm0+ODfw8eGJ1KEsA/AB8+RORYEf9qWJCzxMZ0Ubalhn/tSjI0KVLlxSUaWS4MIPLDP6Ed66L1a9PPRTiNwBb9h3Sh1anKZvwbMcWgVC9SOz5tWfDflBFqKEe+ChlkD0Ix/pY2fdotatWoZYC8mzDu6paVEnaQbdPOrligORp9MCWWIdCdK5cDkHWq4oWUfSfewYfPCMXlHiirWlWhcokAQIBkchs8Rxx8DaKwuCH8P1Po04tMdfLuzPYiaRs89K8AofkfWQUq/PEBNaDbQTuPJhFAAAAwM6hABq+aagQ+/olOIaSQKkeNzBBCjKNdvAMpo/3E8oojlh7RQcQUDWKpCJAg8eS+k2JT0SPbaLQoMFz++WX/IaIS8vGw5SCMrhwOQZIKk2oQ0uwJhnxDyLcdRjAEDUsoaWrJw36bwZBgRqAMsiwXqsYgAHyZ0aIXDCoBrRhvTAiPhfohLyEY3gyvgb7Aq0vPkRRIyA60ErHImjsNCswgJR7bCDILD3ogQuksglKhhDCTyijIcollonKaKmqHYND4Bw0DcuEsM9B2iAUNKgyZoZwNJ+psEoPkuygaQz/iQNde0erT146ksei1fwAJVqNa1pQor4RO0IWcvRhylCGipoB0hikaREgqTD3NMMh/AvknGEM6CYTMhYBrjCpP/zHEoFLh3cEYcbfs5B9ggAlG20qFTOiYWpXlSAJkDT5Y/yIbtQIJWNn4tAmVfwhg6It/AhAAYYn0HPgfFhjiBuSEaHiGN0c8unaGHKbiTSKjlIkwGG6nmCKYd4NxtdGDPOUjGALLCYRLUtGoApgMmpqhEz5mlnDUIVxd1MjMKp2E6h3OBO8ujDPemmubtC7toYW86ZqjuWRogZcWAlt7AAJOQMGYHRgqOSHiNGtFW+ISi0yzTrIt5240ukQDmCECoW6qQCTk4xkBfAkEXnjRKFWSfSd/NUKJqtiMOcO4rWqSHVDIaY014IBDF1VOgOMf1sl+veHXUfta9htlqCSRtHmZoIUJePGDiDOeiUWNRYkC8iiJNIP1woSujZVBmnnObP+EUams4h8DqjBm5t/GTWiEUGuOlwpJqABGkoXGHzoFg/4g90uTr9XbqNADCWQXXwLwRYA33gjkPbW701s2EjsBtseAt7lVsFjwBF6MoCkRLN4EN/Oji9htCbB6EIM8lQs+/IwPXfKS9SaHhiFU4RbBMAZVplCvUaFhBuMjnwEkcQtJpC8ho8IeMCTipW5NYQaUABdDJjEFaQFgB3ILxBhc95cWrYYQuUJYAg9YRY/EBRDHQhgvlOa8fwxxIVqYAvLCpS4V7EZdkDJGFWpGM1K9sQqTq0IKyFAIMBSiCtcaQWPelRB4kYpoyADDIAtBBc0V7hYLkYQhmqKZmxnyH47/gIyPpNIUAExBbjsIhC908Q8qXoQLDAlleBgwSiueEpWobME/DvGpf6hsbv8oASwXYjKiSAUpAgLXtaYQiCo8I5HBuJnQ4ni+QiDjCv9QRBN+qZk/MoQKrfrHEJrwjz7c4g/ag+YQcNiHhTDSjYbEVySdpy0WzKApNWtKIMChkgbkRCQImA+v/kFPGv0pJjWxSJxSWcWZNIJsQVlIhnjDgi5q4R9AmAJCTdaZKVAISmv8hzuYSSU5UoGbkvCmNW9hgybcIhA1G5VBsDe5G9bQIH3ogyTIYJBoDo2bErnFLVoqzDfywhDfW9keW/jMQDyDnQtBE7JmwYBUtmYinyzL/8TIhoeC9bMsc1kILx6oBjBmRg0qsASnZmaQDEUNUrkwyDOq8NFbNEESVThfRm+x0ZS2taIMKaYkuFnNlF6zCUMgKQ+H8IdqhsCafQhBN8bwiybwsFWFowIVXBkgdRrij8IcQxzcaZA18LNrnEDLAVCjVKiOpFYLs8gCTVMPT6aSF5YYgQqsCq4MJXIEJtubQW45gjWSIyF5+AcUdgsFUBikEC1NyEdDkMgqxPG4lUvBDWf6j0QGdqU35CEZ0ndWW/zDFk0Y7Bj+4QzDAiOaBkgBD6nAx8wgrUtB+EcnghCLQKAgLp79B2kNsgiRjAMtpowJZ22SgAKOBA8V++xFqP/GEfOIxAT/wOdGAApVP3CBF62UWkIW8ItnCMWN5k2IJEdQBdx6JB8SIYM7wjAGtz7Xm934RzcIu4AYuPUfdEjIPBjCCIM4YQHMNGQhePiP8hpkCmowFxUsYQBetGIH1ZBb60BSi04uxKgWoYVseKXfmPiAvyPpAp3e1B2EDZW+ftFiKkMJYdV+imYtBYcvnhE+pHk1jJg0RiDcsWKPANYgCxiDLuwAjlHU2R196EYfxjCGGMSAz3awAw8UYZB4SGQVFiHDYYdQaRz+GHCNMQR4xQU+YzzjGQE0SLFEYt+EXON1avFBS7aMFtfR7h/12cNfTNDqk8DzJAL+xzGSOmD/02SkzLy4EgSFuVhIgiMGY6hCIOoFyR5lpgdR+AcPJgIKGyckmY02CBwesegFbGIBLo4BOJj8j0CxwiCdHIVBIv2PRzPEtP4IRx8WwNJJ/yN9aAhCtnaAtMVmwADOnhwwYrGLJ3sE3b5WeO2Qwut/xBcqtl44fv5BFi5wYR9U1ReROU6FKhTCIGOoqPX+0QqG/KYHShiJM+yQcEXboZMH11FCZi6SwjITmzw25L7v5+MgiNfHhuRFBtCwAwBsEte0tQk3UEMWg0R54l0j9T9wgQGSDMSyKwoWrD3CJtS0wJQXNyoBiGYJqmaAF+37xxiKWzkfG6QTrkyVMTg5koQv/yRQErFDzUXCAx5sgrt/uAJ5g7BH9lIhBRlIQftSYKpcNGYSSIQvWqQxZdM43Z7t0exqIhF1jVjmYJ0Xidf/sQS5owXqBpEnULH6jxmcz9kz/YNeg0CFIARhpJEZwTMKG6yXb4IMYOhxNF2agiwYIOALcbZCaiHfXoWoPfo0zWB6VRHSJwQ5B1SYR0Tf4JN4DDyeGBdk1BCMIADDEgYhgS1CgNYhtA/x+/jxP8TY4XEt4E4qTrcuQkAGvS7k9jIgA3rMpRKiE/jlH7xgClAgDoDFCnwl9TwvWErA61Qm+xQu6RICoOTjGsYMEh6hI/4D9SRiADwhCnpAM9SgFc5vIf+Q4R/8yoaGIODkgR+GgCl2QM6eAcZC4uAOrix0ARz+AAxw6B9qzwAU7yIWSzieRwVGpxaeyGCc7h8yAvokUDUcoNUkjiMCDC0QauKQCioiQCP0yxPIgVOSMCEKIa3wzQCCy4a8pJfqxTTyriUWwAn8LyGOMAMkQr3Ua7GKMBg4AyE2qRaQwguBDCSMaqisUIDS4R8c4BETQgs1YslQST8kYg3CrEyCJSOMCvp0ilwmQr0MYgiOyQVTwHDI4awwAHuWzQfLoolGQheagBGoK3v+IQNYMCGWzyBG8QAJpIhUYAeA4KpI4u4YERkVzg8uUSI0UTYSjCO+oyN0QKwmghf/e9HH9CULKMwduuEXwIHcDAXdYkAcCgHo9hCSrhEbe9FcHqMcqkEZWIC1DpEkFjEZrQgSbyQW75EkaiICE0IVNIIAF4KHgEG91O4fwCEVWIHa+E5XFE8XOcL2dtExYmUSVIAFlkAL1MBkZCvq1GItREEE+DFY9pEkbUKe/kEQ0KFj/IIVXhEtHBIkCvJ8QIIKDODtGIk6ykEFZMAKrEAL6FECQfIke8V1nK8oPeIMKbIsZHI+/s+lcNIjhi/ovIQ6sCUHNpKMPAIpb0QtQHI8SqMrTQMMkxKVDgwk8qL8DIIX/iH98rAPpfIiYHLa3mQU1REkOsEQ1OB5cmCW1CAo/7MiJcwSPDIwLBxua56KMDcCLTsCnjiFD9JPMt1yIaRyFA1iICcCF+gwRWrP525SJCYy6NApVh5AAkYgK4EgK5xxMUtj6tCC60RCGk1DqrYmaixiLGPC1BjCF4xBrFoh/RZrMoPz7T4C5tKtI46R6mLuTUQzh7qnHPwSMEOrNbHmL25TIojyIwRsWFqCBUivNk/LItygTm7jAivmKbDzH0xrPzgg8xKCKWYg/figSgJOreSyCDEzX/azOMuCFTjzTkaxFb6EOkaABaZAAALA+6pzNaaOlkgCExIKCjfCCTyCO23C68qAIVjCJP+BPMMDMzDmEgxiQjViRDUUPDJPFf98oTv4QD4tIYZ+7vb0s8jeUjX+E1CCZXIC4VoUkAUSdDAZVIB0bSG6QC1EISGoYSGkzSIqES1eAJ44dMw6AhoNAh46ogo1AjNEj0RLdCJ8QUQQgAIS4gMeD1/2KBcMgIfwswil0kbxsiWorZOoLUc3QirhNCbu1DMrshy8QBlUYBfSYA2A5T2FtCWm9IvEQj0XohRCwknDQkJqpwgsYL5aolGR9CQKlSEqIhg6IT47Afn4Mz/1pQoIgAIooAkoAAOaAAMA6wb+4QbEQRz+wQXxrCXoUkX+0DGeZxIsgAbSoC40IWy2ZtZUgy02Yqh2AjwmATEN9SSAYCsRhlNaoRX/TK8VjCwP9zMIxAEDfmAN7ECKpuEd/kEKhOEf6GELTtUM/gIqJeEyZeNdce9d0GAKqiHy/ocWXMdGuIAsZkFTReTupE9F7PFgEKEWUC08+MBOUAMHstQmJhRhfeUN/qEHLKEVomOPiixU9TNfqmABpuER6sEeNIIe1vW6SKIPhIshXpUMcEBWRQQ04ccoMAEEaAAONMFGslQKkOUCWlI1NCDLhGohmHEjYjMsCmUjGnUhrs8gyjIpiUIFikAokFYijLY93kCsZsD0RqATbJRj0yoTQPAfmqEC5kMP9IAeakBb0aIgRfEW03G9pIZM3gAPPIEIVikhikpZD8bLyuJY/50VGaUFWcB0rHKhBD4lGNKvLZFvTU9oAR7hHZpBIughPWBhPNSUMucDkvhFbgDgGGIhEVoAbxOCqUCCDciTYDliWAF3JPJxImazn/5VJAS312gH/PYjEPJCqt7sFhdCHJpgAcb1JOwKKihXuN71Nnjo9tJxQOVmErzgQf9hAFoCFD+CPf7hBDzPatHiSu/R1FIyJrwUJe6EUnuAEs7JCpAGIROicDAACSSXRtQ2W5G3PV5qUewVE54gS7OXdUfiNf9iNxNCaSeiWEujSXq2f1uiMS1ArEZgLvigLf8hgsdrCChAGPTgXOdDGMr2H8a0OS8TDYRpCqjmATDhBVCAY//Cgw0SGC1MbsBMYYXbw2QitD2EwgK8jA/CcyGWawjEwYN1hQhhNugmx4e84HlzIII5Ar/C4iwmrlj+dzUmUSKaZCEelSE2jyMQGDz+sT00UTtLYy9gwiBGgBJ4QSpJQCLwzyBIwyCE9zQ42CCQYAtkg00v4ucWq1WCoXmVZBJKoAMQJSHU5C+w+DbENoZb8wKY1iJMIYA/pD061CJMGD8+VCy+WDVQoAo4ZQSszC/W9bMID49FiEC8wAtUgBc+ABLKDZVoYCGauHaatSwoNSG+4A2UoQBS75A1woW1uCg14G8ZlE4N5fzw+KWyZRJihVNSeQ1SWID6IpedtW/FAnb/Iw4uUvciFvYiLtAiLHkjWABFY+IHRqQ0pChYkO8mba+E+KUcQicKxHANLE9IrTjqCNksA4A6y4ICZakMENioZNcmUpkh7GFcxxWOfaWObQIngSHgcM9+d4AqVCAQTkcVUCBaizJCaXgjoPg2COgeMfovDFMsFLk93sEeQPARCpoRkW95o4kKrLIcgCAKhuUaGtPz2OKXNYJJD6iAB2xiWyKnFS6cJcKNZeMcuktXVDrgoikI/KYqvKAHwHSmyabdYuKmLWJRWViAIDksFHl0P4KNxfAk5fKgNaJ9kE+ll7cTWoEvfyYQ4KlEl9jXqvoi5BmrueYOekIkuqBKR+Kb/+taLP5v8cw6qRfLHUcgCgDaIJAUv+R6p2mErg3mnoOFA57Z88QYJFzhH6R4I5ZyNgGZJHbWGf6C2oLZVxgvJPaQ8QLbAO543zhjCqLgBNIAD1pEFDRALRabISqhABAh61SEZRCGdidCikEPNbDYFMjGo20CEFhTIl7hHzDVI5AKDFf3HwVZI0iDjWWDtBdC1NoDKj0CtQN7vALOAPwGB3vgVwMMAUpBA8bhWFdtIQrgAg6hzjpCq9HisWUHBzCauFWDDY77gPL7I5Z7PhhgAhiAixMiHCRCDLE7AmIArGWjuxdiu3tlD6dp8VT7JvdtZjwhey+hCBDAAdrbB3wZH//+YYm5gBJaIBfOwJpLA64XjgtoGEhG1L8TwgUa+WCSm2vAcAAm4MChTgT/4QrWbY0X4sErDMnRIrsTosItYh0YAhvmo30u3CAU7/0ar/EMwBL4RQ3a2SC+gAscQBTY25dXbRw0IAG4oBVmIBbIAUD9WjaE0q8bYUENIrKhgool4D5mYQK44MCn8A4o1QIIHQdsQI0nYmdlY9BO1iBsQBHAQJkWgh3AQ6/0yso1YggUD8tV2wDodQaMARzS4BK+AAHSQRRqO9VF4RW2oQUudgbKYAaeIRxjA1go29cEALO2t58i1dfu/B/y3C+A3MBLaQIG3QJeINlBQAhwIBxIY9H//yHCUaPSJ0LbFuITEsII0iPTLwLTOV0AM7x9OkENGmPUAwAAuOAVHOAVXmEOmIESXNRFY2EGSmDWuxtXAbx2erojtIbXQ+KJKlrORQLYxaKxS882/BzQDfzYC13ZXwAEamELkkmNd7bJRYQU/uETPmHbDWLbM/4v1hcXRx68syADTL7TFy/9YiEXMMATYgGCKeHx0GkG6j3WZ8BFcb4K3qMudqEYBuy3LSJdEuLfQUJ8B34kAIpLF6Lo/4FIN2IJOuDPD3zqjx0EQOCGb7gW4gAHnIC7yHU+2OETJF3jsz0hwEDsN54U1l42vvsitvHKTR7lEy/DDWAE9NiVXAuC/2q+5uW95luBEHThHpBeI1z3H1rk6AlfJERvQf6h6UFiLqjewAHd6r8g60GAbo1hqvcDG7DBGbDBFiTdCBQhtHEB9M3eCD5BEcYAGx7hG06j2ydiD7fx5LPA9lF+0xePSyiBerzKqmYgfW+eD1rBEKAjF/TjxRU/oZZf+csisqf3Iojg6TmCCicfyO+gCIoABL4ABHbg6mPhEEgAeOcDctdYEbTtD1r/EbDhG7pB0t+n0UKANEgkPGZ/5G2/9lE+3FOgXACi0z81A62oGXHQyowZsQwZSPGPD59EhP7tEvAvo8aNHDt6/AgypMiRJEHuKIkyo4WMRVKOBOFy5IWYNP9r2vT4IKOXjBh1kKxG8oKEf1z+TWAwgQsXZocsVHuzw0JUFT1UFB110+W7f1s1PvrWraO/R/++fXOmKOOftGH9ZdU4JAtJeR2zyMuCNy/eDFkypEBjyBKfg4QNjhgxw1AKXhka87HEawQmmCA5cFr0tiabzDTfvOEMmiOQ0BovzOR4krTqmMt07vwXCcUAzk80Iv03QOmsXLwpuYnVo8eIJ7kSrcpYYfVHso8eYbsX4w8YkNi+xQjHTlEIbMpBypX7r9DGLEfImy+ft7GhYJRaIbYyAv6IwClSDGk8JEWnFJRyfB7JwT+mZBRgdxpxktFmBo4EAGUL1vSFckzAkBH/Jg9eyFFOXmw4CUa4aaQAR6GkdBoDRmXExQBsHBfLPzME00pvuXSSCwkbSYFhRls5100IK4zBwyNueYWNHdVtxR023D0IXiHg/SPXEf/Ic0SVVFapVxB8UMJLMGgEQ4UlKTyUQgb3NZaBAbzwwod/qYGEYI4ebebCPwlg+N9/co70mkd6gvbmTV2Q5EdGk2j0lHJeLDNJowI0ogQC/6Ay6T8KhEjTEh0hkNQQ2jDDBS+W8GaIIbHMyMsVHkWQ0QLdcdfVP81tBKuszC1JFi4LZpCReHhpJGWUVQ5LHpb/pGDIDLzsc+yx+dWHJl+LtZBLCf8EStIiBe7Z0QE5Osit/0YAuBSgZSnV9k8BG/1p06AxAbVaOf8cMwkAHUZyBgKhoIJpiKjMEZK1IU2QEQNKEZHLNswMsQ2vU/7DDy8JrxouR7NypdGQF9IF5cMcbzRsyEeIEax4bAZGl1/5+YXmfSnsU0lE13q0ww49eDSgnIuwwUmdGo0TGifbVozSoSlhtsgsI6Gb0Wkzy2k0JvCq9sAyVS/jBQCRRLqvAvx+jSlHQFlQgrql/TOURhJYoALbnr3BRcMZZSDPNinE0gkveXTEakYRuDqSrqqR9Q5ZGS+4zZMeicERySQjI2VGkWfRSTCPQYlfy2buM0QuGbXyz2dv1lxzwQJuoCDRmKm2Ov/RKRndkQAebmQKB6mPxIdq7rruUUsPXJ01vvqCDfY/nmgkOwDjWvtEAU4L7EcHfhDhxyFEHNKD8oEws03i/OQikSUfseqM64/gsqTgGsWqHF0fc4TMRoyL0YYYyNAvBskapQljMIztEy2GIQMURWHCP9xTOtIp0DZcYAMbhvYgE3VEFP8AWkmw5REOSDAkBuQdRxqRkUhwJndn82B3VAAEICwDa1rL1766hooXIiAKARBADQWgPBXA4DQXcF5t/MAFBggxKUo5hAow8QUcTiFUfGhFKzrhsJTEoG8LMtw/NJYjuihuI/fLyP2+iL/61e9+YpALLwzRxBlQgRfyyMD/NrQBijy8AgEFeMIFmDACqCiwZlOYiMR4MQttmChAbtiT7bKCQZKAgDICM6EjV+OGk4yrO6nRwj8eELw6DA+GXgsFAgIRgFDKDocqKMEF7GiaU0qgA0IMIgIWkRsiREGJkElWK2aABl64JAY0seJbfNmd95UEGfz4BzLagMxjtsGYZGxjENAYjBm0ghLbWAUd5pCOWVxABk+QwQiUMYUdqGAEsaDEYnhBo0QwgxmcUNo/JPVIkezAQk8byQ4CoZGVZEQG8dQIIGDzlpMw7R9P2AG7HtSSB0lABVPQUAv15YIXxjCiA3hBDW8oO7I9wY4clYEEEhHEVhqMC0a0wJr4/zADlCYGIr3yyAJwhKOs8ACLIxnLP3AxpCVxi3EZ4WnkNBI/ZbaBH8gs6jGPADmSZWBUTUzjNHlBiYxAlRJcOoSoysSPfVhCMessygb7aU+NqKAmYwXrwMwaExwmlDQqKGsmEeCCiEZ0oqgYACHeYMNRCsACLOADE055ylio4BCuZAACkKKUf1ACpSqdQRB02THxuCQCUqBiZmyaEWCi1SMQaENnP+vZZLZhZFUyUy7ag4Z/BOOAEuFDJ/ZDtyPwY7b/AIanQgrBzYaEnroFDcFcAgMmDLS3KInQRvT5j9GE0BNwlWsonCsOQhCBAMYwxhsAIABMsKCbG91oCQabm/8gBnIbXHCiE9MYDEtEMSu8jAHgbuLLd7CPuPD7R2g/e0xkkFFk6OELr9bLD9nyAxnbGAIgcxHEbaCIKP9o0WYTWRLk0hclRakISFbiYN4FYE8P0Bpz4/rcEMe1olHIBTknkog1tYAXK14TL0CqjRhv48VUfW0r0GiITgyhLpKtyRRBU76bPmg6LolfSZaZEc9CAALI6OxQAwy58kSOSv+oEjHb0OQAi2MbiQhELIrCCU5AQxtsKMo/JKwcM6MkThP+CA5IA8+P4MEioTPr7JRTVo3A1QMg5jOfxaGDSBgjWdJ0bSeoClVRKZoSieASVWvcCUM8lmM75sgW2/wWCIz/RL9AdYmmM6LpT9tXjPkDlqmbDAoSgAIUmj6CPPhRtyEYmAthng1nJvmGXTxS1/9YpFj39IEczRnCe4pCuJSxkTq5wAPPXbYH5ICCSBTjGbmQpjnXZIlsLxqqlqBEt79tiX1QyS6YXtAmFmfMjxzTvh0xckxEXWWQ8NSYTIYAUfkBgQwAQxzaIIqa53wTCwE8JBIsVMXIyU/lyCE0BMiIrUGi6zm/gQURgUFtMlzumEzBuItYtsf5vAgPEAAPjSiGoC3BHroQs8oNywAXMsCYM4mhmEQtda/W+w+c0/e9FwoqkpNcElGHOtSgZrcX4z1aIzd56aAVgzjc+I8hqBk0/8YFycM9mPCMk4TYGnnBhTbMrar/wwMZ8QDIRb6LRgACEI2Igjg+wDCk0tsjNjK6MZFMHpL02IML+EWrNsJL17nb3f+AN0oMn+QjYNm+9V7yktvQPW3MJimgMYZLrh6TOU/SJo1EiQg0cr2Gl1vsHLE15rX+DwtnZHUeQIDIL6H2RjQiEoGogjiGADlOj2SZhM/Id1D/jyBn5gbD7PTRNYL4m0hJ8UHFr+O3EQoF2+YjXzhoSMjOrc2DBAUGOgSGvMEZC+gaXMDfCIUy0oMckGTksZd9IwIgDvv8NCXI/Afj9t7bBfRN+B15aU1WoCoh4W5IxmT/EIDJxxEIaIAb8f9z6QZ0jmdvyPAp4rBgH5FrLoEg2icShfJmFYNmI3EnI0GBGUEEGyF6NhEFxhYTd5ARscCCXBdPJQgSeLALczZnH9gRbNY6sAcIcbB2bCcAgdA9srWAqgJvdecRDagRHyNMbUZF/CcSQsA7AQgS+pVfyNR4Q2AM4mBwIqGBnHE8LQiCI5gZAEd+oTFnNPAPl4AIHAF+JmR9vHMzedYRC7cRVechLJh5GeGDPtgIOIQHxoBv+nUcH4F48xYeltYxH4EE3cFzNRFTWidqvVd4TeZZhHgF+BQIz5ARYcgtlteJbzFnoAgSf3KGxHWKPCEuyIN+b6F6cuJ1GmGHH3FnMQH/e3wYB3HwhwCACQCwA8bADKtQiJzFgLwXbx9xaRgSDuMTfCFhWeVXX5WIZZ5FAhbGfWfmESiAAl9IGrOYI7zWa+FCfCCxYWCHEsFWEQEwcBwBcHdwMyL4DxQog6sBQpyBEZP0jv/AgnQYEv/0D3HAEbxYBJNRe9sACqsAb59Wdz9nZPPnMVukYCSgKkjQiDmCFdDoEaAAEkjoZAMGAatQBdzYHQBXgxj5daHhC/+wjmYlQlkxSbwGgwFnAUWAXYFAANZEB8MYgAvpgHXxD9LXEZX2D4/YT0S5WUj4D8MIgfr1kVWQkiUhg+ZYE+Oykh8xj2GzGrqmhhpRlRUjlSBx/wmkBxJPyRH5qIIucZYjMY8h0ZJZwWs0mBFnmZYc8WbeGBLKEyFz5nUEQABygAAJMAd0IBLzdhct5SSFsA2SpWB78w8VSVySABJVoBGMYBMKGBMkgJkkAAGauZmgkAu81pYkQZY2MWeXoJL91JWuE5oGYmxziSFYkBIosJUicY0CgAcB4Aup6BHjCBL1yBO2uRFhOIJ9KQ44sA0isAo2AgHbkHvxVghDIB6FQAY4EA7hsAWZsAnCsAAVMAr9AFY1oBGuoBGS5ZAZQYUcoYQpgZQZoZElkWqZeQWqBgHPcF0c8ZXdUYujyRFkGBIKFgVvkJL6SROmCRKewI8m2XUocf+CWQGbJeF1cyagHpGaCwJwFiaDDTdnuxAIUUAIBCBr3XMF20AGGJAEFXAOzdAMzXgOGZGi6+AK3tlPsPAPg4AD5yk58sNFQMduQaURNlp0N2EjqrZqmLkKeZAH22AMgaAC+FSO/3CfmzUi5MiKHhKhCJoVl/ACZ6ARrukRC5oRsVgSDfcBGPAPz0CgJXGmLrELKbgaUnkJZ1ARFKARorcLNECgGQoCgYACOoAFW+ARUJgE4OkEHeGYLgGeoDEITuCjHRE5lNiZdKBqqiKppDGkq0YHeRAPCeABnPgPgWABXmeOIrSa5VaSrPkPxgaOImFhr/gRZLoRACkngaClGrH/YRFqYQ0npyCBfSERBmkKcRlRCxkxoRuBEU96E75JqwClEbDJqv9gp2vopP+gjbsAAihAAfQQiRuxov9AD/8go//ADm8ho4f6D4dKrhnxrSMho4PKEQ65eBqBZZ21oyTAD7dADlu2anlwHETXEYWIhDayaqn2DySQB6BAB3QwD3nweT+JAA2KjQDXlqO6EbkaElw6YcN6qjQRbBnxAc36EdywIFW6EbqGmySxsXIisSLhqyJhlx3hj1/pm2Hgif+QqzRAA7XgC7gZANp4BijwAi9AAK7gp/+QohtRtP+wAh7RDwtLEzKarv9QAclBtOewDjVQA0/bEStgBoUQP8OC/3TpNlrwY2+OFz8QAApksAs7iwKeQAA4MAShcAVGeqnX9A9xFLB7I5gHe036mgcKEKXdYZor21siayBkio4oAavKEQnGOrIl4arhaKWZMbMZAZs2Wws3ewlqqwQg8LMU4ApmsAJIcLRQGxZJG57U4ApOaxPdeg4nmhE/8BHNIAzdirQdMQjUEAYoUAWrcAWQY3+/a3c/53yb2WSaJg6BsAtKgAKBAAJn8AIgUKe6W5zFOQQ4UJwEQAjHswspuY7smo2RSxrBKricEQb/MKshIQ0xAQcgYQ0bUY8pmxFK8A+EyxEOG46SuSDFsFnZEBLB6r85SwM+67MvQAHicAM3gP8DmlC0zZAE6AoLVlsDqDsIG5G0WLsRsPDASaAHrku0KVG0tLsRg+AKyhsAtVcIV7AKNEeJhZdk9Va89Ra32lAFy0vDSoAHePCmz4ABWLDDFEAIFBCGacqpHdgd/ssRKXm+KaG/9csRNxBnu9q/GhG4N6GbKCGze4KsJSG/WXGN3REJ/mgTVWwT8NsRbdgR+ASmGYEDriAM/yAFFVADmUAPFaAHNZC6gToIE3zBe1wDwqAHzZgZsAu13OqtnysENFDCz0AIz2B7VzAHeXAFBQh08XNfm+l4mqmZ14QDnGoRF3EG9ku5dbAR9KsaASonXiqaGhGsVGy+NFG+/1C+olz/MeubEWD8IOJpVj5xE2mQBh/xT6pQEsUQrLqGTxmBAXJKATfgCjWAIyj6Dw28An+8oilax7CQtBO8At3QrX98tOcAhUQryDVRPsKwAq4gCIi8tjuMBWGAAVVgnCLwyMkZP6oSVCRQvPaMyfEZn6sACttwvDm7EesMy1iwxcA6v5zsElmcGbj8DwwdGg4dEk/JuCqrEQUNfLTsEbNZEoLAEWPgrLpME/ybEombcbRwxBo9sa7gCn9cASugxx2MHP8wzVC7DtuaETatHM7QDOcgBeC5AhigA8WgA4IQBkXNzsl8wAhMBoqKnHybnMlpyRKZz/nMz6/gAVVA1LCcEaK8/8W1sMQoTRKpihJn+qST+xFLfBNE3BH6+5TBGgDjmyMcLRJybUKrPBJ0XRN4jSFd7KxvYcsZkQrA7BJ8TQGFXdiukLQrILUZUT6jOxLfrBotnQTkLAggRNSCUAd1EAZYEA7J7Nk34NkY4Au+sAtnQA5YgAXiYMAM0z3Vq9qF/QxK4AtKIMscYdEksYyhEaoeQbEggdYeUduuI9jgCxJqqNHD/RFS2B3WYMvt6xItadcazdc3QdJwkIsdcdxm7BFhUNjH7ArUcK7N6NgfMdPjHRLCB9k3fbTlkwThMMeZgAGrzNF1QNQYQACG7Qqe69lbcLO14N8569W1EAC1cAldLP+baujfUvjKmv0W000Tdm0TxWDSIFEHQ/tIDi4S1lmoF9LLLgF+ZDmb6DASmnATs6ndtfwPgMDcGXENudjhKGENxfDbNpsZL64RaUDLIr4RiKDdIj7hGmGzOnDUn6vBHVE+ybHYG1E+wmfTNm3eGlEBRRvlHOHYQQbHil0B5KyGUqjcRG3YK2DYhr0F/i3h1kALwozmOOsTIN3Fyq2lSYwIIq0R5CAS2Tq/Y/wPwuzcLtG+El7RbwHhGiHnLqEKqaAR2pgRGM4RqOwSJE0Sa7AGGL0Rkt4AH4EItXACGpHpyI0hCl0Sjajca43dD/LXHWHowHq5J0ADOkADGPBmIPz/FjitEeWDI+lNEiu6rQ0cFnrQ0ucM0rdNpscs7PxNC8WeDbTg37VAC8f+CzQeuUkb7CUR6iTuEmpomiXHv77p6SIBzILNa8a9GiQuBBHg6I8OB3Bg45D+D2vA7Zlx4jXhj/9U6jXh3Kqgv++uHGlw6h4BsoGtCtaACJegA4igCSrNrbCe5CiR8ByB3rMOEuZ9tC29AuuAHDWAAZnOEdQe7Y/rrMVOCyAk4Y1AC6qA7B9h0iCdEaF+5hph5tQuEoiwlYH+EXZOEiFQu6abEqFeEyDk3BMOQn6n8yOhCjqeERjvdy6B8Rrh8v9wbhmBCC8u6SCh7hzB7iHRyy+uCpyO/xJBf/QhQfMbIe+ZkQ3Z8O+D3hEWbuE2sb7lnhFpAJC6EAeqkA2IoAqZYAauAMJNvycrapQjIQyu0A1SWwENnAkZgfIakfaw7A5xjg6qAEIibw3/zuMngOlgDRJJn+0/LhJqiO8cYfndMfeHDxKJHxLIKtKi/xH7LqC/oPkhAQmEmvL/wOX/gPocUekkcfvsXum3rxFVD5DcINiq8IwawQoZEVNSEFN+Z+i00PWk8eJVHxIYDwhaLxKF/w+CoAlmzPYi0eH7zhHogA5x4A7s4ASZcKjd2sYaQfELstgLD8gfMfg4/w/rQM4rcAKOGfQZEd6pcA0A8c9atmy0AP1DSP/rxL9ftH4h+vVPFUKKFHUgRFRR4xaNHStC6hjnmsaF/2j8AwQozr9GKDtyRIjBI0taLRtNvDhTJ0JNJXVmo4hk50qEunYe7Qjy3wmlSGc2+AfV6VSEcOKkQQgplUZuOiMglEIx4r+vVM3+g3PW2sSOYztu0lj2H1akaZGm0QUnBg4nTtf9+3vWo9CZFagaDlyh26Aa/4QhXLeuG7VMTjVVVHUQnSp0FLOxVfVV7tHRLgXr7PoPpNyy10YifH0aEC1rp207TbUVIdGmFWlN3XpKNdh/YcMSR0j3tmA4cFhRVKU7Ly7lS8nO1L18pt2Ka/5Fo9jbrBCKjysKTS24elH/vGu+NWH3h2I3j3/Xwf2HJLD2neYpGu4IQMgGWeGfCtap4LFNknDlH5g00uQx/zoCpLNsYvsHEVVA+u2fa3TzaSe2guIPIdEQ+Qokooi6Dah/XLQNiYwq0i29g3BbKT3+eECIx3981Amcqko8S7mR6DIKF51OQCQ7jQSkyBmPdIujMyF3koo7J4FDSEDCEFpgOe/GRAutNWJwQhGE5PunsjaJ1Gi/jiacKsEuhUkinCQ82rPBx0oT7LWJovsnFUK3Kg2SEyJisTyEvtRoxkH/ieNKijDEqKLXDroRToQWCnEnQCnqrLNUZnSKm+dQEs9Tin7oiDtXO8qSolWTY08j/5CaahSsZo46BRJLOzVLGoROSaWsOHTrzKkwT4NKKoS802iNNRpYoS9bKgrHLChnFUyYbuijyL4khFnBlQKFUVQwFpc9KrstTUNoxKOA1OlWjxptFtypINUotn47CnWu7xDSd96OhHoMYKpWTYvaqPzVCLyK7PhHl2iiMWorj2HV6NYInPn1145S4TECXcBpVN+jpoEjDayw2ooolnUSriIppdRoYMGsbYAHG8DQyIwQ/iG3oj0pSqIGRczoZpO/vqVYp3WECWxP/5LoJt0VanBFCoWRunmlzlblYStLO8I3LoqOmxKknKuOlz+qZ+qsV0BTwxhjSrOiqG3tTkFWI/9Z6dZJGjiURCsaOLYC0setsJIGF8ZNrgjkY4uqCB2idEnDYqfAM4qb9ZDSvCKXzYr22gYWcILNf2x5eiqu2emFFEbYsWWdBfYLTI/HlvZIasgE00Mn/EJwIple2DHDFXrAfgzz01bSRV9jw/sHZCCJPW3tioxCaqVep1p9bBN3Eo8bHXfice4hD7Z1qgWMe9Yplw9HPNZ/7GgORWCWsH/cqiuiA9xOlGQXlumCKNyR2FGotTrbsOI55HNKtP7hnQZgi2gIscUfnjYup9SgG07oRS8okoy+UMR4gcEPQiaUhKvJaSr02EkSVsCIf7CDFKTIhzqo8Y8kZMIV6/hBq6brogujGMso5EvFc1IBsmCpRn3FQoqSTvEcVmDQI4LbiRe7lwqQpM4j1utIGrgRh+dcZXXyu9j/ZsI4qozKf/+gY//MEsGOsEIaz/EbAv8Bx3+8o34a+VzEyGSWAJ7FH5sr0bWwYQNF9OEfIdiWGQr0pqTxiYiZ6IYtwJCMfHSEFJ/4hCLCEcPjHW8FKxDeP1iJFB0Sb0+bCEcyoEBKhDAieiJYQRJ0OAhheGwqV8ILHDCGC+dEgxVY0YXkClUoMFIsDXaYWTRmZjCKbG8m8mOF+eZFSLd1xJmnQxg6t3IrWU2jI0oyljd34o+AAAAh+QQFCgD/ACwAAAAA9AEZAUAI/wD/CRxIsKDBgwgTFoxEMADBBrQU/mvwbxqcggAEFgOUZqBDiSBDihRI8ZLAY8sExhnJsqXLlzATqlMQc1FMhRJc+rk5coBAnyy1CAQAiCTPowcREPyFtClMiiAZ3pP4baJVmHgGSvtnL2GPozCMQn3pwanZpwntnF0bkkWJfznZyp3rdCzduwiPCZwksKPANSIB/6u3pqhCwQktCPxy887AaRVZhp0b6iBFu3gLEiHyjzNngzqU/OuhItCOKeWqAag2CcCkav8wKfu34x+If4Ge5eLCJZSCVwn+zSE4IrPx48iTr5XRVG/KlAUxK58ukLnZyiOnEkwkkLtAQkcrP/+RMFtg+X+wBaZHul7hbC9ecvB5YtDNcur484OMAJLNXE4wcaOQXnJZV4B+LwkFEnYIIYbgQQAIIAAAx2DCEoH/YCiRMtAhlFEPfjD4jwsG1dNSGQ+mCNMGSPH3AnUkprjSXej808g/3gxkjYrq/EPTXRn9w8I/U/wzWzkKeYFeOUAUyZKFFubnBhf+xRiNiWZJgZQDKhpH0SNXPSjATwTRVJmIA+3yTw4KuqRCS9qFSdCBAtF51I2CgdklcucVVM4IfBhCRSxICvRAocsgWs5zhYJ0qKGFHgpdOUiWg0mjAlU6UErpBSlQAAEIUIVSqcil1D8MpBpSKf+wWgqrxlX/8s8FA9HAFioSXSbnnrz+E0dVY61xzUB2tgQYZE59luJkBU1QEAqxFMfSFCxYQsk/DxDUp0iFYppQo8o8oEw5RRbZp7gDbZsQAFH0OlAXDyUX51EsgqSru4EhZedF0iUknX1HaShQjRIt48g/MsiKX5w0xFXQTgJBjAtM5ajBRw/kqlsOugI5eeijU2Q7BaC5EGnQA1OoIC3KgaDRyj9oABPLP+SOoAbKIxgiKBrSEqSpt9Htii9CHJgiEAcCnZKf0WcBxt8/bw4tdUwfGYXYjgrJ4ZQJAnEdEgos7NFCIom00MIsLXCRth/iBEJItEvY/KaTBtH9Zw5GYqt3tjT//8PHFIAHg4Yh/4wQzEBV/APMP8YMVLMhwRgSSCA9/0MFGkNI0kQTtxwOs+CWG1CIQGAsroZAjkwxQyzmFpSypwdV9Q/sPCk2lylI2zR1rxPsZPvuKqrFK1RrKDHkPyj+c3YiLJwOdUHSxvLWQCMURzf1ucyA2hQz39JHH1QYbrlAktjyzy0FNZH4FJEXhEYVVQxBBucCed+EJAYIVAUwQyhyC/ro68M/+tCEIfxDcFRIQQqoQDjizEAgQSDI4daAGbwBjyDMaEo7/rHBf2jggnPx2lH09JL2gHBPzmIAqibAhX/MggvXwk0sCCfAgVBOUP8wxAM7JpARNG4T3QBDMv9CgotHYIMHPFjAAmKwgO+F4HtjWAA4BDIxVggkHP+AgkjAoD9J/IMM/yhE/nIYCCIFgwoJhNkBPfePKigBMP0qCGNc8ju5IO2EeBRJ8uqYx4MwBS9MEMhX6KLCFqJqJ847IzAiOBBbhIAgwKCCAVJggAYWaWZT48E/FCGJIURSIFRYHCgPgoZyjSENFGxALWrTR/34IDO0owuX8vMmK/SqATMyyJjuMsuR7EEhH4hW4SwBjDFCUCCiRKZACjGEWyRxFAP8xwKUsIB/TCwkVrzLxMAhCRJcIXNU+EcGjJmQcFJiBuQazS++UYs3WVALtoyXSF7Ax1aOpIP2FIgoYOX/LgfNRYWtDGRCCqkEIRCiBzOwBDkVdxBGDsShBrnmnsLJE0OMYHss4EPcrBDPgRBMIf5xCZpEYop6sUWLPMFnPllyPMb4ZWiiaEkcC1IbIPzDpgjpiipFMo6B8NMlTCMIFlKBgpIZwACWeOAYw1lMiSTzmCtViCjRoIaQjeAJZbDCCHIQJaHt7kUEudhdVNorgblLoCDMSdRw+g9A+LNLIOhBFWZQguK04qgJMcAQyOEPXJyCFf44hZboQY8aFBYWFDCDU/rxDyeQgQw4gCwZhiAOceAnCMEYQTlUwIcdBAAca6CgifzgB0PuTmH6mWlCqga8eoJQdwNRmkgAUIR//0wvj7GgxAjewgdLpKAgv/2HXjFQAYHQw7jT0QM9XEEGSXgxOfkLLkMPOIIdjMAXaRCEHzowAWcZBFkgGYZAbuMSk0bVJUtQiAjM0kuFvKiMCAnpIgDEElqZhVXtjckvBxI1mFwPPz04RC5GMIMZSDIDVzhLDP6RiaNoUjnSlS5BDDhdCe6gGiPghR+6S5ATRFV2pTqviI/zBoHU5qMhKUCxjDPIgdx2IEE9y4OTINsRw4TCBzEEGoKBmgf0IAq26q+NY3Ib1x7HrAMd8glNwM8NvvIlvFByZnAsECojJQhYFlQneDwCFfjhFf945ZMJgtr8HMCebQrJ72oLkzKUwf++AnkBWKeDyd0NayQijClC5iiQGIYEPPD9B3gO4gzqLDghY/hHov/xSBsgZwhZkEgGQHLUIBgAy5a2RDDUMAM+aEO8/ziAD7rgB0pc4AwULAg4RlGFHuxGPzEasZClzBNMdPUsNxpJAn76vOkUOj+k+EQ3umELdhiBi13axj8ifQSBTLogWTBgCoag10la+6hJ/YcloswHv8WCD3xoxQzE3QpwdzoWuU0brVeakS8Y2SAQY+lZRHgU+7bLJUrKG3IYMIECFAEERXjDDkCwAxXAIBet2AYJVuCUvibkEf4QCJhwgY1HPCIE7ADDJxTRjX+8gyDv8IcznGGHiFvTLPL/OEizU86SZjd72VnIQMwzMG0FpiADvOAZJXiRAl7sYx/yyEIhskD0I8ij521jZUHMu+6hxbIp9/6HrEo2pHevlG8hIdHTZxUSFajAAj2wwBfwAIIvvAEPFmDBBZ7whAtwIR55+AcShmbygXxcLpEeiBiQIoYjHEHozy6IJ1uBBl7wQx5H4McqqhCINzi+jHx0gSnYAFsLWN0pnLgjcgJtG56sGCmsBYlSSiYS+pylpyoqjlCwHhKHgAohB8rFiwfSwgH44QVnt4AfVpGBoRP9HywH/ir+AU2zbKLpEGCJGNogEL/LI+i+J3oW/N73I2RgH7ywFiU6QYVOWIIK1gIG/zCmzYwMiCMW4shFGRvfdL9J7SPxXmErd4kgoDSCFpEIQP6/wAIWxEIGT8AET8ACKuAGCMAFB8gACGh7L1B2ZRchFsAHvMALCIcGM5ALKSAPynYQ1bRu/CAGyIAQIdgSJHAQyZd8AsF8/wCCA/FyArF3BAEBMjiDM8gPQ7AN2kBfSHF5BAFQANYUn/cSDGEcJfYPZzBk03M8CFEWBbEjN1ILAmABQLBVLOAGzMAFE7gPlAQM2WctXkgJ25cLhqBQ+zAQMScQG5hyedd+c1GCCOGGB6GCCsEI/0ACEGCHdiiDq6B4vJB+4uAHhFBiRfh/TcccLPAVTwcvPhITiOASW/8REmoCEoMUiSHxAXMWEsqiHDPjGEpoEDahFBRQC75CEIbxD0VQWxYQBW8AAC9ABFywCqtghwghh3KYEC74D/nwD8c3Hfzxa+cFCgbhhigYgyh4h8aIh8iwD1zACeJAAIeABf9QhNEIE5TYEvDAhjdxiSPhCf/wDP9wbyYREzjQErZSDAKRa320SwSAECiwC7uAAvEzfAVRCGVBAcJQASPXDMX1D+egB/+wDgWxizHBWC1RAwQBCwdxBS4XRiExgv9QiwVRgiSQD3RAB6AQdwIBjBkZEhj5D8D4kSQQkngIAasgg8hwhyQgDiAQANwIQtA4HXyWEAQwaBgwHYiwEkX/gY4sYStrUZP/4JP/YI4hkSNNoY0DMY5RIRBDSBCigRA0EI4JQQH/cAPU0GAC0QwCoQcGCRIIyRP+aBDNgJUKgZD9EAqF4Hf88JAhSALpcAWhcAV5EJfJl2DDOBASGZIQwAgiCQoimQckwJfpMA+r0IwUQAAUQAHt6Au+EAC+sAsE4AT/wIT/oBRlMY7kxXkeERI6AJWZsY4FAVsh4QsvwZNmUQcI4ZlNAQg7gjUtkWiBRgOI4GEIsQX/gAV1cIQ80QhCKTW6YBCA0AilWIojgQIDgZsE4QpJIBDOUAHF5QorcA4DsY/MKQxJsJUK4YtmkQmu4ApbQJpYIJVNQAGF/7AKeSACcSkCOIADN3ADWPCUirmYiumOKBAIVfAM8EMBhBAGgZCYtUkI+DkQL4kUomgQkaADvUIN2Agnf5EGF+ESAyqbdwFNf8QWmkAQtfALohgRMpIQKGCgFLACrkANrkAPXykQ0HkQwjAQKToSJ8qiA9GiBMFw57ACGACh/1Ch/7AFDKcQA1oQtSCaOkCaBKGhgjAQgmCcA6GhUSkQtFkQEEoL6DgsBloQOCoRTToQg0AdtTCgPdoSqkAQQlpNnFkQNzAQHnYCESCbU9orkFAQvTkQkGCjHagfT0MXdyYSDdoX2TQQvRli6KAK6BACTuAKVtlxBiGQMIGoBVGiAP8pEAC5j/9YEJD6DxWwAuHQYCvaDWagCVKwpglhnQihpAfRpgchBCBhlXiRCtegCoAgqiPxpV86F3/6p9kQE9dAqgbRiC8BCbh6Xr1KEFIgBZMKEqkQqy2RTXuKFBVgozwRWqHVDezwBwNhA04QDtbJcKA6EJvQqF0iDI0qDCmanP8AooNQoa6ABL8qEquKDiH2Dw+WGTHQpkozRQpxChHQriohEG8qIHeKFGIZEnPqEhBap/9gRcIDE1U6EmAyDVUBXtRRFbJDRP+gJ9GQrAPxA1SEDQaxFdJgRdnksCzBCmnwpmeRBmlwsH+hENhgA4owECFgPmawowRhqApBbAT/kYsF0QuMgEUJsQ5JAJDUeRCKqqL/sJ0pmqLrUAOuMERDJBBm4Ar9QKj/kAT0AKIpyh8R8GAYqxAWiwt2oAvRMBCs8GC44A8ea7FyYUVhiwtrMA1rEA15WhD+sLUS8Yj/ICAS1RJ0+w9ha012+w+p8LcE4Q+pwAOnELgG8Q1h27F5CxLNsLe8EiddGjRQ0bcCUQQCo5MD4Q1QqSvkZRCXELcJehAj1SsdkhDptRbJ02tHoTX4olrUIZuHNhKyoBD95Rh3AUcD8VYiwRcFwbtwcRCfexBvxWbfNRLW4RQkgisKAbvUgZowAQhwECcRWxBz8CMIwgJxsUuWu1LCKRAo/7tuydsUD3C68gST//ABuGuUFxQKzHsUh3AX3jFrIqEk9vsP+aYQ1eAFSJIysTAk1WNbozvAQ5ZLCrF1o5gcwEvAIsFK5hsS6eG7CKEMSBYTXvAahVMA3uFdDNwlp9LBBCEgCVHBIDEvsIcwKgIwEiEUaXYXmUgQxUCUA8Es7DEJmDAJjQI0+XsSA0HCEsF6BMEXFjAAIVUibPHBo4uvxkIQV4ofwys1ceK8TtGbX6If9DYXTwc0PlMcVFcNfYIhYHwQ0MEhA+EFfbIaABAhuyAhjBkA5lgLDBEJteB6xfB6ohl6YxIFA0Bf0SDFLuGDqCISH6QcZfYPWQGyeKErfv+cR7VaEN17E/eyFqG3lH1kQSHxBsIUEuFCLjqzODmsxXdhU+ehLiMBAHdAAJCwwAMRBd0Gwq58QZEcCDKgYkOTrl2iCsbQX6SMEN12OkA8EpggALswCeFCJLqsbxxjJCjzJ4FSOemiOjPzXxJxCeF7HE9sEIpoFMDzAS9Rxf8gBaSHH24QkyLxCJOLF9+7FpzrL/9gwkOhIhF7Ai0mEOEMoL8wp9JsEKJMM2rgzAqxzCPQCjxGM+ITDFVgWYZiJKgBKANtXYMjEO+jQIAzArkQC5NDOAf2VAjhJBdMvP/wDbpAQreFVu4SYwgSa1PTAQVhvK+8UsRjoMwRSLnQz2v/UtM9RBytYMkIwVYEQTdFUgX/Y0YNpD8U9Q+20LJDUEYPkDMEgQZN3Ukty0mcpEadEAT7kzmMltVDkFkjczgpwEZ6g1MsUA1TgJlW0Zs6fUE6GBN6RlbIodIScc1nMRwqYkLs2NIt4SyzwAuxoAYq4DwD8UfSYmB84M//MDNNABOk8EVUYAxVgEZogEZD0D/0IxACNApjEAL3IwnIQAp0+A9XsNj/wAjJQNrdYAfkMBApEGloZFEdw9QGwAuPbQnFAQ4UYSImgsgiAZoFwYM8wQFrfRRn5tYtERxs8QYWML74wR+zVxAvlU8Eexc0fBCzBGYxgTRssA1XuA+TTRCF/wCZWV0FhyNKDBQIdONDC1C95WxNuuC1msQKEyNRurCnrECyIWGoCyZAYMBJFMU+4ZQ/TUVh4VMOO0ALqXZCPog0SLw7iywXcA3XUnMwycHBI0HJL7G6TXFbB0LhHDAL/3AIsWBBraBQyrQ4o0MQziU6zjVZucBjBo0+PGHf/yDjN8Gy/0BhQZBA24BXCaE9mxUIqdAA7izhGREAz60Q4MW+eL07+7TkUoYAdUAO0TICxLRQlIZHwEBzL0EFQfA3lFLWu6ACHWXTMRF1Z7EIugPIDT4dqpwccYHAUqPETu4SqT0DeGUJFaZMev4PELXnBXtyNhZBrQA4RVIGGpUDp//D0wqxAcGNEBtE3HOeGXYtEnL+D2Hh2yER3f/wAjSOFxhQY/3CVh9hU6TeIFYxzyAxyE5BCF/qarFtUQb2Wzg2RotzVMXUVPkD4MJ1E715sL1pRZ1OF7m+637OM4DjNyXAVQGADm1u0gIRvwJxZtMhKzG0B3XGK65bEJqbH9J4EJg+YuklFEGSE4rerwMhwvmhBF8aAOSQPQSWUFGm2gRxVOKwBafgDyd6XAYhs2uh7wLhCgVh5XeBaTy2A5ODSg0wDUUK4RTuEvXMEixSxJEuF/8FZ3Rh8TyRXwrR6GyYC51QV52mQAfBPzeQCT6brS3NSBSlWSqQCx9QBYTAzVL/GQaZAQ1smBUvQdciUVu6XRB3oHQIcYmsVEf+wdsI8TJ08Qoa/xL7JRAOUx0gFAiKYQziMAQn/g/OMLsD8TQLRqqaPhcfxx/DiiBWBkFoBDPaw79fkQpY0ko1thZyPfEdvMM+BRPNHRMRALkGofdRVfY3/vciQW0FQVGXw0BUwNUj8wTMAGrAg7spAudIwdIjUQIYTityZuYHwXQjwQQW1O0EYQoA5SzKzSsiTPcHwSr4kBCAIbpMgOFO8fVyf+PRlhCWxuW2j2WDXj3ikA4eFGoC4QATUAlPsAANgBmA8Q1roERsMWaxnxBj3vwJkc4i1nE8OxeifRzS9WxreGM3/35tlWYAxXT4FA0NPqAB5v8KHVAJuRAFcaALv4AB4l1g/hcLLZBBHN9HqH4QFpIVkA8Q/wQOJCjQwT8LBRUOZLDQ4UOIESVOpFjR4sUACyf9i/TQxEBMCL9ILLGQy4B/X0AMBPFG4ZiLMR8+wkaz26d/RozYqvdo4KZ/OAcqWvBOpsxtAwsNlDexUIYMKaKmMDDEANUUhv61ojSjlVc+rcIGM2RpX4Z9lgxR4qXCmMBFR2WGlFvX7l28C02xuZhrYKV/Pe4e/HfwY17ECxUkFohA4IQBBL7s+vKm8hcVMHJdqJRozkAk/xbI9Ce39D+fAnEVXC3Q52nGBbMoPGKxtv+YI0cyPJ2dYQjBIbwMxTIgj1kWeVmOFDqSpRCXRFMCvZnicC+n2A/5Yueb3fv3gtmy+wU/UcC/83RjT1H2b9kyxAUEyoDIqwcvfszk8ZN3hd//Vf6TSIryCrStNruQUaiNf3ITI4ssdssgQgoz0I2XTqiwhJdcBNvhnx2k2yEWLjhhgJO4BuKCFy4oESeWDxnjwsCIAimIPpmI6IBGHnssrzqJXMABhQAiKSaSAAIQ4AsYYHiCiQueeOIfFf5h4MoruTjJjxcse2OXNwQAQZwAt9mPlyoMoSIFOiSZyJl/4IzAR8TyaJBOgcRQ8E6BZkOQIAbbEFRQZNooVM//MgD/xiwY/wEhRjwjrUu+7xoRiACFUJJrpX9ekIswSR/KIaWIsBuIlkhSDQAPFVRgQYZZONhnH2aY0eZWXLVhZhteWqCEklYMGUusVjqRSqCl/mkqO2fmtCgGOEM1EBkICBJjoT1JAIUOUPLhNinHBOIiFpccFajcirAYCN1MCQpX2oIAKA+QgTISyNKFuLFoF3jv4vQoFmA4it5/xPuiCAtU6MFVC6pgZh8ESaj2n4kLHejamPoIrV+OeWTwH1ImlnhkEiReBYIjeBFHyyimewOPjgXrmKAbCPogtmkEumQimCtCwSIL3npoMTp7duiZf87A69F/KSBADnFukCMpbgWa//gfQ//BGKJCul6KhH+2EAiomcGDgAQ6wKZRZIrPdnvksxXATg7wfLlLHbyU/oeGgX5GDNOyB6LBU0+P+kBdwwcq5t7AFRLPIgoI4nchpZWggJoaKhjoHIo2XsiMgmARaBCFRBfdLhEubhACUEpGBpk/BdqTIAhqr9btf8BWWyA6VqniGRy2WWWVV+hIOw+1W89dIFD+yQOU53shAfnn015lG3EsKEbJABYviAAiFrK7cYiMdsh8ifSeCHHEFwLcLkC88WagjhaqXyEdFOLbIQwKqiM2fJEvIteISC0kArp/3IAamdDcP4RRA3oIQ3MVEIZdnNGMgvxAJkkYCOnMUP8FMq3iCoW4wuv2BAoReAABHgjeELYxhEKsIg+rsFpBSlYy5LUuh9qa3vTyEA864OAftTDgQjzwD2ooBATq+4e9GCOHdx0xL+8yECL61qm7CGIi+ZvZL2gUwHup4l4EOwoR8QeRmkXOIgRLg0Dyx0UhEMSKViziP7hYh/f9wxWuqIErVvAPDAqwgivQRDiUUMcwQCRyajzBP3xRC1oQsRhmrIUOUGBJN6KABrXwRf4SGbaBKGF8ABRNRGgxxH94Ty51ZEwdWXkUJSStPFqMyT0GAoe6WDEmcdRfx+h1SkDQYn+C+0cm6qKLuqBjiDSgwQl0oMAV0CMTFawINb+jh4H/YFMg2hQILMKxjn9UIAkrEIQuNeGjcwqElwIR4ym3SJBGxoRA5NvZP2hhDXcKZHH5jMko44lKiZziHzwYqAAdEgeKNMNZMfgHJP7xT5mQsSI8cGhBUoGnNdxyINEQiDRwkQY7rGETTmDHP8Bgg2IShIOJIZtDsAlOgTQwIg0UxjqSIIyVDmSPrvgHEuYpl4uqwlkEUYUXK0qQn8pFl//wokWGqoo4pEKZA4FEUh0ixotYdSDphAgBlQmIoQpkNBexIj/vcgpWNE4aBLEDRwsCCYEuJK0D+UEg/xFWgiA0L9FIhb6yg9C5DiSj/xgsQaaxhjU0oBtOQKlA/vAHJ4Au/6f/qIFKBeKEZBTkD2NbiDUd+FmBeDYm9LAsTP8xij8ORATU6MY/6LECV1RAgzEBh0IEOtfA/mO2AomrgU6B1lOsxg7/SAMr2vgPZMoFockdCEEh4gwpaFUgrPBrRTSIUFyiZq1HcYbnyGdLxkGkAQJx60A2cpSL+qie/3jAP+RVWIOCZ348ckFsSnIRP1ikFEehW10c8Y9GwJdjHCBIPf6B1YqAaiEJiW9BjkGQ8QokwhaZL0HKaw+B3K8gObvLhGOCopiga0r/wJFcUDGRREREwA9Zr0BWjCcDEwQEEhDIfQsyEoV8ciD9i2+V/pFdggy2v+H7TmsabJfxelghRf+SCCCS/A8lDwQIERHAetea0W+Ux8BPjkl9BXLiI0PkxWGGCAts/I8Hb5TMMqmHMdcsExrfITYAOI9gBxLliCAUAPIqiIHHrBCYFa4gjchZRtcQhzoPRGCGnQiOFp0YMD8Ezz06BKUoMoIR/CPTFkDB5AayC1/EIbkZDcdnBHKYBLxZ1auWlqYk4oWCTHjC53GinR/CZ/AcVyAM7oHMCMsxLzskyhcQSIrBcwiFjFgh1bgIswUC62p4QRkWYIEbBsAMTgRCAOpRiKVjwwJFs1rc4lbGMtoLYSinO1IfKLGBZNBuxEQaL0RmDAumDOuB4NvZsdl3SMqtDBXwgQ8lGNX/QLztajw1ZNwLF+CkCZJoPJVXIFMtT2E9XRF5R8rU/4hCtJ8dk31XBN8XgfUU+ECJf8inAMj+jjJwzPBVH1XVSs4yjnH9jzgMlsMKkWh2gEwjOFw8zI/+R3sogomNTCLa1TjvQtJMkHLkBT5eUEEsjC0QL4PZVDIpA8x9lKIvq1qK3tnZMW6eFzfYrCAT+MeOvF4e883i43eZBCaOEfWFjHzk2cF7NT6g8H/U1wUuAPvb4TVciJgCMUuF+csrAnGL0NgibQSEeKzRRI7AAcOSyniPWIB3izx9IeXwAt6fvnfGlP4fUQc9QQBws8APnjGpMTxjFK94YavbIj7mEZhD/yGRKf/33AtZgyp0aY3LW0SvEVF2Xuz159oPpPkPYT18/qGGTPM+InQWQPcFcPaIJB3p7WG6exRSjgfDehkh4bZAovAPTow9xohZAL0vIoqBdCH6AsG9Qrh8kSiAN+d7iN+TiP+KiSLwDm9jDIfbv4FoPYhQk0xTP/ODD+sbiAssiHKwPggUCKO7wAcDgGrYM4EQAH4RgACwm8WpNYFAqDRIAziIgzMIl7iCPpmgohlZM12LlroAPIloQJgjIAj7uXixCCD0hH+IJbyoH/BywBIMhFjItIooh1gwhCAwhCloLwvMjuEjCApchnLzwAx0CKNzPRAgghtIL4hwqOkDD//8y4uksAvSckI6oTgJ+4f/kYjCOo86Wz7EoCUn/JeIwKX3a48uHIgyfMARyAUqAJH2SkQDwbsHKIdDrIsdCAO88joCo0PDU0O5GK/5y6jCWUCOsb+OyS+BwCU4IAcWAJJKVAhlaK9YsIR/yMKj6Duje8WFyMUpqA4pfMSia69yoEQHpD0fSSIDebLNWzUbXAiZqws8I8WjAL+eU4gMvDofaUKBaKp/IDqIgBSBaC9dZK9A4INGqURIhMWiK4f2GMYeiAUVwLuoi0VKBJJafIApmAFDQAMqmIEOLIcRCIaFeEV8a7875JHDSIz+wwuiKRAgVAjGiw1jYxeKuATJ+4f/iyyQ+ZuZBzjASNHGcNsK+fCEevqpGPAEKSSIKbPHhVCDGUhJiKgOSiyHfFSDmQRIPviHTrg+gSBGfJyCWJiBLKRJgdQKQzAEYPDHfOQDmxyBnFwTKgiGB0jHDpSInRsIATwKv9k/U6SIZgwyK3q/F2AB8uBE8lGyCiMIbAyVESgBFngCSmgBh0ABJRwINYCI9pgyZehFiZDEKRgBQwiGEQBIshCIRlSIHXDKXDAGbQuEYNhJgaiCKviNYJgCsjAETAsGKkCDf5CEJpCEKoDJgWBJ9ioHFRAlX/AFFEhNfrER5CoIJoiv2/uHwrMI8SBCs/yH/pKJh4y+CBuvrwQP/wUrs3+4AErANClEzhxATuxbTuyrRYXQS0Usgbv8hylrr16sjiqozHzUCs6MzH/IAIG4BU0TiF68zH8QTK2oAoFAA0kYAs+UBDdpz4GgAvi0hX8IAUkwAIH4L6D8B/IQvmUDkRghB4jouk3xDrn7h9kkr9zMC7abAFQUOvF60Ikwq1DhssIqga6bBT+IhbusziqpTvP8hzOrRRKVsnwUSkWUzD5oAk2DSSqoin+AUYGwhVuogl4EzIWggiqoCkkgzz4IgSZQBILgxyEgg4J40SHAzBHIkBQAhlYoUegUCMEkCPLEpQnTPvJZ0O/QAI7JKDuMDVQMnDG1UMRgooLYh/9DGIG//AcroJKBWBmBGNFYyAXXLAiTk8yBcIKheE/wVIg+GNQmCAZDNUx+5EdggE8bzc9BHYNbkM/JHAJFaIJbIE8hDYExWAC7OczfEAhDsBFHUIPu1En2zNF/qK2BuEo0VYh2+Id2eFXyacPs0L9QEaOqDLJ/2MpWlYsZYbt94IUn8LGAq5l/yNMRoAIq0AqFgMJ/cIdGdR4+iQgbuIVgAIZFfc8msNEhPS2B0AXE4x2KkASksc9P/YdltZFejAWBSIFgQANmPdZfSKx/YFWZqE0ewVeZ8AGBkFVZlYnhvIvjqjN2/Yc98A5bDRwNQwweI7OElAkGmIBZ4IIM4AX/TQuGGQgChWAogXBMw6QCTCuIWBgDO7CDBRgFgThXSfsHO8AFO+ABHliAGHCuf2AFXHAuO0grI7OIdQoKEgAGUD1WKUyBFHCIQECHBmiAZRQILbgLWvAULrXQVHPCE/A1lXTA4JQJgSkxDCWIhD0KtstBLsivfPwHY4BMhZjP+gzMgVCBESCEf+DYidjZ7xgump0TMnhPoI1KgRSIpogKoAVVfzxWHkCsgtACLSg4uRA071jIN+vNVRPE6LPB5NM1mXgl8OACceDJ9GxEjf0H/nSIGd2GDDAANMg0oGRPAcouRfiDTz3MlO1RnbTJagiEWkisKPPIXv2O/3u87OgA/2RjsMBp2rKph4cciaiVCNGsCygZiFmIFS7wQQKAR4FoBUsIXY0FBknA1mk9AkDtg4Gwgd8xhlvwhZkNnBDozN/QWCqIEP78XIKAXcEcxilQAjhoAFUi3hTFzd19u0RYy4Eohf2CF8Wdmd5chimbCASlEwTAgmdATg0xgNCFiMB1EwOtrQUYK+bimOEajSEo3fCMCUMg1fYKBF8ohqjVXYuQ3Pg6AIJwYe/I2u+YsiXIyoMQhVJ4w/79ByqKvgmYEXKIwhmwBGCY4OhTW9i1CGCgAmA43V4sh0DoARZYgiWwgji1zsBhgxQxBR+0CxiWiS9WsR0W2F/jkYYlsyyziP9UeAZjGOLA/Yc3vgg/HQhWYIUNhrlGFMxeBAI+KIMqtoLEnYgNCLzumIh/hYYxjpQvSMeIwIFMRMxELpABFjOI2MRNJK5AyAU+uN5/gNc3/uSBgF+JUNW5za34CoKXpMl/4IOXtIIcIN6K4KKyAQyBKMtIrohxGAiQLIgEtK9QESg8s8emA8eI+IZasFqJmGSZcFwCS6tYoAQq4JCAtISi/QdaFIgJnmBRDmW7CNfpes2ysYT5nYIcuIASWIIcCAl62eUwGzFKyIWCjeQi6GUBis03AwJ8ts4E9sPAyeQMyIUSyDRDqGbQXQhgEAdJiBqERmhJIANxIAOIFgeVpQj/uoWIKtheaTEEoayOJ8iBHQgAQDDcgojesrGle8CF9zNgdZutMoUIyLvlxNCxujiPVsFIiQAjaVEBeH7Jf5gBCYYIA6iCeaoHzuEm7xAGPaCHpNYDpq6BLYCtOOwRjQ0CqgbZXmSBXci5xBqslo6UYJuIg5UWyH0I9JmZjIS5qIaIErjigpC8s46IJQiVHsiFXBiBGehkXiDodh2IISAAJOgt1+KROfwHbFoBG5hoH/lctQiGHQiEQACHBrgHQfCDDpiAH44JGAZTudiADXBcSUkHVmPBiiA2A5nSr7sIcPMvaXm/QGABSyiBuy4BYzHigVhUcXAzmMZmguiEjTaG/zNQgjOogzrAApmuCDDdOosYZE586Zd2CGVOjL0kiAsgNvlIXoLw7Iuw7osIWIg444eANxzJSokQXoJoB3wojyoBAWMAaLseYr0miDxIHYGIVgPRhN2aGdr+h3idgkkYAV7oFT+wbIgI41VLLYvgVzppyOwgTYLQboHQ4n8o5IggtrAmM7cjsbzIZc3+DuElhLoOhlxAhitYCI6NALmVibE6CtPqmPdG14EwhE6ozI0YgRaQS0/M7VXj7Io4UTLjAjmbCMxFDOsbQ5l45IHYRORGDGdBAmEwCh5pqY65CoIAhiA4TDRAA+6cBAu4gwXAJRaOZE6JEbkMnC6GCFvObf+2I4i0U4gmRL27eIIFLohLzouZPfEFmCwakbgGY98rf8kdYEdzdPDdldw075EiSOD+/dpQ8YnmFggcgIfnxpMTt1AajV1LjwjEnvLPVdYrv3I3/cshkIV/8IENN6g87Rjwswt6fgiEewjSFogXIG+IkHCL+BBidogLF6DqWjUjjw2aDZVMxwsqqPIq30xUdtMROAQ6mIdRb/bHoAQ3OIGkXYgsmycMoO+j+FeBKHULXXWKYLCsFEuISHKKiE1b79iFq0aHeIUBjnSCGCWJILA5l3WJ6HUcv3TRNYCqrnJLiMK25IV40IAD0GwH8ANKeAIdmHaBaEIeIAcCGAJtkBT/5R63HMwLDo3NnEwMFZiSC5BGr1N3xHj1vJAuiXByuRAKUiCFXhgIUiCIli+QYJeJFFBZCZbgGQ0CfbeEl/RvOhj4A/CBV/CDSriAM7jfwYqAZyCEEQhKS7AVmEuIWzcQC0hARJcLto6Nt65VAcJpiKB3s3z5XviEl1d5Gon5glgWhxBPbLaKmpfgIjaAnSSRdHiFV5ihGqeERMiFKoiFoCwDr5gBPsiFfZA7Wl+1Dzn1hzDIey8QZ3O8vPAeN78IxZ+IMiefaXiEEACDnPiEP7CD0nAGGygpgfgEMOgGbIANOpkNglD9f2B91ZcKor2KmqcKA8jJTkC5nv6KKdV9/8APhv/WaF6gBD6YkUWY+MUPFRzzermgZQuPicgvj4iNWDcoAhBQCXNxlX84BEYIB4HwLoiyCH8w+bn9hm/oBs03AjAIgSwzeWwIB5xQhBXABh7AhrtgfYqwf2WRiAmBipkHiBQpDAhMQSXYjE58+Mzg0+ofpRQZ5GWouC9XrkQ9/nH8t4jjBo5s/HQsafIkypQqV7Js6fIlzJgvQbDk1JGFzJwqu3CEp/NnTC9AWXZAOaFAERBf3nxRaoFFrgsdhSApKUXnO5iP/HHciqsjtn9fv77z9yir2KEp5XVke3LbP7cn5R0xWfffkUL/smTgm0GiSQPBglliKy/LkSyHE//LSzEkV6B/FkqaUju0suXMmjfDZMNxEWaYlf6NKDk5p4PUDjizbqkA5ZtqK5+U9MPrkKVDh1Qw7Y3naYELlS4w+7ei44LWQMP+ewT2X1auylfy+5k3S6EsWYZ0TMExRSc0neTRLZS4ED9msXb8Y3+6IxtTnv/Nmq5yERub9vdvBnAyAH8SsMcfSgJw9AZ/D/yj4E+yxcQAF3JIEMUIgbzxBgBvjMCHIZbksg8oUHRUwT8kEggUWvvdhVIb/7QhBkvItFEXjYlpl8Veew3xF1+WGJJLCvxYkoMK/7zhXnscTcAJA5x8tMgiHPyjzA4qxGKMha19NN+JJ51GU5cr+Yf/kjc1wZTLP1LlwkeYJhm433vKeLGMZk9IVUkJKHGBwAQdvACCMYUUsk0G22SxjTx6mdTEdF+lFVOKbf5T3UnIvCTjSWK0eARd2PX1aXbaidEjFYZQwgtEucRiSCy8MAANR8wwwwUXvPiYi4c7DCippHnyxwCvwa70wRddSlDkS6HgAEIAkQTgjQABCIAJDBwxwdEFOP3DALDA/sOnHy/0BoAxCKyCI3YcbbNNqRDAFME/MQg7lBC8QuAuRy1uiteN/R5xhBhHIMMPMmJYys8R/MijMML8iMGPwpZUYauu8+r0nsX8EVESAhnDtLGkEvwzhUsuDIBCJI1E4qyzX7BQ/4IMMjwxMwsqfEArAwhAiMAAfqigFIa7CACAlbFss48lrRjCh3cqXcWRMx4rJw+MrZGQkqWTdlR1SUe00QYEyIQ9Nthiy3jEPuJsw4UbmsmGoNQWd8zRAKwxMEHdcbMEYJjamhQKSjf8k/LKKwcAQA8SsADDzE+MgEkstCLAxc5c+NFDICPEkos4trbCUCvBoGHJPh0pilJy/0Stt2VZu6h31jC2QQIodIACyiokuIsMCaus8g9c3poEZk7FqiQ865YVkHxLIID5AkuHuOQT8yd58NFnJ1mjsgAqqDCCBInMUisv5Z9qPi+nUmIJJZ243wr8aBhiQF9xcYRja4xyFP+BM/C65P8/IiCvkqzOY/hayQEPmBIYca0kLerI1e5FAtrlThvaoBUvMEIA6BmpJLRRS93m1pIEdOkJ1aqZTgjQES60BBBvAhDfVFKLkhCPJbuoXktOQwiZRIEjMLjDRlKCAOyhhBaA+EcAdmAB7/VgQ1zYhiW4QKk20EUe+8jAPvbBjIWZRC6ZUs4PmNeNeV3tJS1SoO7SCIFVQIAE/BiCJcQxhAHs4IYniQVLXIBDjqAAJdX6Bx5bQr3XuIQCKWnEm2DCwcwEYhcggNsedfJHtQACQF8oggVeoIIo7OANUdiGNtj4O5NYqpQMjCQqg3XGq6Vxgm1kYwYMIA4uZOn/QEtJ5Uvw0Ef7qNA+rLgER85gw+Et8iQ0iMkdmGdHO3bEGK2hCQAEAAICEEEOclgFHegwSo4osIEuKcQVOrKJf4xBUscRVhmFBbZ/SLCN7tTdEbahrLydhJk5MZAv/iGAXfLHmSw5Jh85A7LWrIEj3ACmS/LZETxwxJ897AgNjgnQf1RBHCl5aDL5w8+WMFQlnuAMQwMAoB1uTA4EuIE4CECIGyAjDxNMCVw64gQcmMEVrljBCjKxhU2YwQmj+Mc4cZiHK+ThH4xwCSleQoJ80GE66eyIu9zZzntpcwCHsCZHBBfMzPgCmAr9SQII6RJIzsuQ1SsmZwD3kon+oxFH/zwJ8RDakkvcsKvB+kBHKGBWFKBgFzS4hABuSAhxiAMHOHBFBSrgjHP84xzNUN28YLESyaaERlmg3e7+4bqObJab91IgBNlpO0HZDhQmKSpHTPuPp54EFLSboCtJgIxVgCIP26jCLiLRkY8OFJf/qCFQNrqSjrKEEBTYocWO2AigyNU+wnVJDBM6nejC5KsoiQIFDLuCZjCWsRxJrE4oy5FBxKQGNVgHR2rwEmqURHb80N0VVpGHVYSTm53lphrzC9sykiCb26BASlN6gyEgQBxk2IYH6mu7eLyCDvF4cDzykIdQyMEN/oyJWX2rEuLK5Lk5wQJHQNylGXYkDSvJ5/8ildCRr7IVJc/QCV6H0mKdALckGc6MiP/x15So+B87vIEZcHDO73bkOCsQ70vIWxL1CsMkBTwJYx+rB2HUAMkcoYYIGPEvgdXFYEeAwHwL4QEEXEEEtiuj2NgJwTbuF7auda1L4UyHV1wBB88Iwz98EQDrxoTDGj7RCZqrGQx0RBAmccU/eqmZ5S43uCzJMYjrYBJC56QY/8iGhi1dkrf+Qwd93ipKhiyFxOpBCkkYxCDWoYd1mPecQ+YIPYRBosdC7R+0towzKpCEGvQDB+TI6xCuQFQIXAEZ8c2DBwyLgyHgAAM0CMAuUPAMcTghnLW99j+unYfa5YEOCZgvfRH/QACVhuG5VZBajnH8Z5T0mCOSZsm7LVZOjpzgJYYGyrut8Q9O/0PTKuOIbjvCDZbUQtMl8TRETWJWRbewEbRICQoQfpKH/0PQJ0H0ChK7jpvq4dYtidqTh0KikJekAisYhHoBGgY8m0RwLv/HDVxxgzDQoBa+sHkxbl4Lm19CBxFHQSBQoAQU1NwXSsAz0kvSYj4DpdHuTolCbQ4UEqsk3TmZIdaZbh+t/hkRHJlxxh5Oi0aoYt85eXg2Hu51lLD8H4a8sVquUZJUqMTTPv+HpPW6AlfggBrqZezIU4Jek5goMwUkeUfIWwFXbMHr9/7HFjqCaBvDnCM574jYizFD/x3QQOLlzCcNlPDux5fE4CyZ/EucjpITpD1M9WJ4sOYNE9TDhPQ6KWhJ4GCHedWrI5HnT+9Rgoha0ILqHhv4SU5gd0HYwAOITsLgB98aEhV+Jd5diSsyoYd/1IACOpihENod9tpLvN4mUb3T1r4SQhvZOF0y/z8obhL4vwQSXx8K/XnVAM7YPyVPC2Cb6IJVpETZld2J2AEccIQuxAHdnYQA/gM6PNwJ/EI4UMOrlZz0tUSTWUYGsgSJNNk5TRlOIULqmMTvvcTDqYL86cTaZQM6uIT4AYX5YdpLUBpKGCB/ZEM24KBLNCDByUQEANC6dcQp7A9LlF3wEQgP8Afyvf9ENPwDHMDBA55EGsRBGugCOjSBCLBDOPxDJpREEnCE9HWgTIxhR0gfiaAXGaZE4ZnckFXAJiSBGRiHFFSFTtDgCnJEHqKExEnNCw7FH0IgvdzgC6JDNuhbSwQiR7CCZvQfR/hg/tlaxjygAA7c7j1hR9yaEGYGD8aENPhgGO1RFK4BNtgAO/yDDfyDGYRDTnHEF36hbwmDGXKEMOzdcbjC/+XEH/rgL3RiR2ziPziiTsRA2aXCAOnEC6YCA3KaFGhCmDijHaYEOqCD3LWED3YEK0zhS0TjBp5EEXKExyXPA2IiRzgKDyzhD5wCD3zjSYTj09gfO5aENqpFHEhKQeH/3kkk4D9ggxMogi3YAkf8gRmYgXqNkUkYpHE4QT70ghOI00t0o0k0GUS2xBr+Qxh2RBg6wSlmXw3sXQTE4z+UoEtMISM+4j/Mo/2lpEn+xDXGBCu05D8gHzC+xDxyBjf8YT2qRARcI0mahDCWHFDgQhGmiD7OSwLunkxIw0miRCiuxDUWpU4gYGb0X0uS4/6txD38QwOEgBMAJEfYgkDOIUyEQEr0QkCGQwh0wzokQVChxFpOJC1eJPaFQxh246415Em0onG4gh0C0EyuRBHiglJ+xQPyQCosIUek41KeCC4IJUekQUmaRGSOZEkyIiv8ZEvkomT+w2S+RE6yRGf+/xl1XSVHTMI/mCZK7B85WgZMDqFrmsQaQKVr+g1MFMVLrIZJJOG84KOwLALy5ASsaMA/+MBrlgRqvkQR/MMxjAlHWAPfUFdxRifzEIEe7ZGf4eY/8MRP5A0LsYS2iAwqMQAH9JZOiIJJDANHIItvoeYxwASdcEQAAIK+8U2j8RtHkOYeeUBJEFFM5MBQqBUq4QBHaMFL8Oc/mMBPLIFJYMxK0BNJ2IfE5c1vrgROqEF7Vo9vSkkkdgSarARxHkBHtINwSgp+qgVzooSHvYRs4lDbSSdH8OZ0+BkQaEaJcsRqTl2X0FN0OoeLqkSNokTAZQxpJmdrYGaPDgWMAulPyP9B8nSUiR2pVpqEPXCEbUIpSgQRLpmmfQ7FmzxpSXyB8Vgp8+Cef55EkKqFgs4LsoSpmJ5Ei7bpSaAVR4gQ62zpSzAofP4D7iWpCoBnTohMmtpHdZ5EPaBSknLEFCSSSQACHOAn7P0DCcGppE4q64yJnVbPJHFGdaICR+gna5RJm7AAC8SCqI5AFBSJCgSCBQRCkZwGCvyCL/iCHECDWP3DHPxDKNggpe5qcQpPt5wIPhbUmxxnyMjpoXYJp2pYIqzEG0yCbBynUKSEfwCAfyiD9xhDLPgBB4QCNNzqR/EquIbrPyxDtHLGyqiFn7YE+gGFDKRS20yH9PwDmqiAMpj/5nG2p39cqHLmRLSWgxrEwpXswBSowT+ka0e0q32UQBlwxIyKq7girGWgJoN0xI8CBXS6hL5KCsS2RrKWRMWmxLLGK2csD0dIwBSU6z8IRTlgbMru60lkbEccZzWUgwowDguURpssrMPuLGu05wNEK4B8LIFklEsc6x517FCIrGZQgmS0rIO4LNRaxnuOa8uixAOwQCswQQ4Y7D/EWGv4Cs9qBoDyB5fERKaehIHmhJdKDXmuBKgOxdmqxIqqxNjqDTRoxMp2xNOmRHsKBczy7UugrElMgjL8K5oUQAHgFclyRhmAbdgCBQN46mbUWJukrXLwm9A+bkfU6rzAxWTk/+0/7C1K/C1MtKfoskS0KkjeekEPSEVHAIvkaq7H6KjsGm1L/OilcgYgnKnspgQ0IAALYMKC6ETf8gfopoQKfNCE/sOgDsWMsqmLcm3vooRNxK6Gbez0Ss17Ds0k0MkyOOtKTEI5eMExeMHKkm5KTO1JCIUKLE9INO9POK6kigx1NSXk0ulr6gdH6K9M2C76bsbG4m9xIm2wCC5MPK0AGIgXVAP4okS0vuecuGdHqK8fcQGsdIQe6ZGuqsQvZO9L4KNp/m9myCmBhEaPLi/rEKhLEDCBWMFDsACxDkV7UnBJCIVsqCz5mi/5Wob5hi5HYMIhcEJ1mvBPYK8H/0MabP8UkZoEEQ+FBeDpEbfER9BuSiDiumouwR5wtJ4uanqvUDhrBHME6E4tDbsEBZdDDHPEQ3nGoNpuScgvYP7DBIStUnaJAU6GEWuYG5tpsBwRIPwbR8xtsHDuiZDM8LbEJHhBIqfEDsesbIzvz3KEnGjGypYrnZzuP6jAxphCdWLAjWbGX2ruHNuHeiaPgjhCR0STb/liSdCnILcJKhDyfrAAm8gE+04JJqdEtBiI8HaEAXPE08pGLtcwR/wsnfztG4DMR2zwZrRtFPOsIzQsSkxDR+xSSHmmUf7E4m7GrbLOyubtCHQoseorA3PEMUzCtFKrSYxvSsgGtaqygSiqSeT/62kOLkdE0xcEcUc4CmeYX3fGRCl4DBSrxSizhg+qQB63xgbAr8cEwGeyxDZnRhrgY+aWxLK6qII8wMSu7xTEQjB0Qi7sCkeobzWEcQ+XBOger0kEM7UmsLSIVCQUg1vt2xHV41tlQyPQoNkBQjEQwCLYRGsGC3Y+c3SqcExIM0w8dEt8QELfXtiq9EqsSqkY8kgXc0dM7EbDREYP78RiwiRgAjmXxLRyRAKfHyDEQRygAAHwr3L8s0yUQkDPCx40oWYwNC4lkgC3hFFL6kSD68Uqw1WnxAgYwj9QQRZvNBlP8EtgNVcHthgvwzevhPqCdTksZ0moABVPBwqjREDH/3WYuO5CfaYzqsVHNHHGtANQ1G1MbOkjQA9troRI8YcO7LG47gLOukS0TsEMFHYwmGa5/vJQlPGCQDZH6HDKQvVLAECHskShPpRrMilRS+fFUmxKBBHRrgRtu6ZSV+k0N0JkHPJJKAhgl0QO8EEQGEIgCMXEAndrAPbK/mxk64RpCkAUYEEodwQr75GUrFB0AwXnyjJL2CkJp8QrRylKvGt/c/dJFIMxlPJJzGhWz0AuBME/gK57C3dmqK9Ga7RKx7dMeNJ9u+Z+97fUUDNr1Gg1ss7iOnP1wMEuUXVKAPbESjhK58QDgDVgj7dKZDWDPADNirFJiPeUdISOu2h2e/8M5TIvr4w4iUvKRf/D8rC4xxTFV6QChSB3R8C4JHPICGA5TPAN6Gb1e1vtFGBrhbs3kT9AFsfEF/zCkcdEZvNqir5ERYvrdd9uiV4D9CDsk/PKXnOElOsNI9abIWd1RyA1orIJyXg5SyxDNTBnOaCQS5RDOWyIIRjCbpeE6k7BQpwEYCO6SRQ4SjS1fWQ3ArB1TGqsdHZABzi4qmdG3A6FKscEKv+Dgv9DoAuLH9y6TnB6lxu6pnfEezOIMiyD6j7AhoT3lPh4hRfzFATCYFx6LFA6s0/BA+j2P6BBMFi7SjA6gf+ZlJh2mJA6dsdE2Q20ZXSA9LZEQc2oFfzDn1//bp1rRiIp9boFqkqsbZCD90loQQnkQDkA+/Dq+IZfe4X7eKXjUS50eZCXQ0cTrI9PQTD8gyEEQ4fEgo+rAB9MQTnsgDEYAhUEARWsxPGaJgrsYXQSkeUeaT2oQpJnjMW5qJ+tW5Lie57QQoqnBKinhMOPTLP/vGMvSMTPwAyogfmWQyDgER9YQiewR8AviMPPQCyURsfPgMVnO2FYQoWXhqLPgCGMDi8AQ9BL8pDHb5OnRAGIO0q8OQ6qwGurRUR78Jk26hpcpYn/QzVO935QD0tsxGu3gEkgXJHDO0rouIzfdkmg+aIvO8EaQmkge6b/gyWkwOJXeKVTfCDM7Ah8/3RHVAEVZMDCc7ohGMMODLYhBAF3SEIwfLfPl4SWIwscVCE46IIqGB1iFqy4dtQnn32wBMAV88ebFNT+zbty8L1LzBATUMLi+kELMH9RHEIgBEIPDOzOW/WDc7vPr+yMWvvKcj/JaPsOBMJui84/DIHYD0jAT8Fg/8Mz7MIuBAJhcwQaoAF3UMEzlEYnkMZgowEVAIQkKrckVfl3EOGUKQcXPjjoRYWKNwB2CRCA8B84jAd7SNj4EWRIkSNJflz0j0JJkbhcqSyJSoFLmTNp1kRox2ZOnTtDAgK5hqdNEzNp/CtDiQ+LGRcuUMrlNFGuWLFyzUg6YmFIZRjL5fiXFf/jlAflduTKJXYEHzTB2G6UhNCRWIXB/hn6N2KEoWBo/lXhO6QJwX98D/KlQqVQoX9DFFWZsdDR11ydPirz8m8HxjdvEAKFExS0Tgxw6tGkFRp1apkyapZW/Rp2bNkYK1WSMEKNmoNavjLsPWKG7o1APpZTUwJkuSm5nlUJpNDuRwMIr4gb8XXHCLoHR/AljIbKkCtkwIAZ0hchFTTAJDX516fPP2Dbp+TlxSfsP4f/dE/K/NG1nRCYDSQGDuJgwKBEIXAk1v6p5KM4GJyQwgqBqjAo5O5TIwfh1AALIRWYuE64g4jjzcTeVNioHGMMIsc57eyiAr0hFDvolluMGeH/gSlmoCy6ugoDZoi34GtCEmAwWo8MSW4J4aA+krSrvlx4SWEG/RDayiEWAvkny4PI+aeBgz7jbYkyMLTppJNSa2dNkspEaJd/XkCtg5o0iZNPlz7rUycuEmFhitwS4o+hJQ79KLKDlJmBBYR6dPG9W4L58qAq3gLpliqMUagVkPz6R5I/EILvj039onGIHE915w9xDAmELgNSoCIYHv/hrb6QyPkFUJ4M/MdN1OBEaMFgEbqEQiL+SUDZjQBQqQedBImWQeQQmiURrFZEqMQReMkvTIRQnKIVYHZ8BqFbAnuGsBTc2yi+HGMc7B8a/aqiiiLnfa+PHJOkQtMhWr3l/1T4xuijCksMoiKDg3J1RA0t6gsSI3LgKPPCBpgdSReVnK2FwGFha8cHbEF6wUHYDoG2C5W9uEykOQ9qWeWcP2qBi1xYMHQjYNjtIasZDCk3rOua+yifg674B4yNbGmiiYD/ydUQNLT2i70hDEIoBHdGiSEGgvpt8h/3Apvalj4WsGOMKoCRe4jpriaR4h/RsGQwQ6ZLY84LS/r4I1M+QgShInQu6didoI0Nk4MgXDw2mkeKAw/KNd95ln/4yK1EkIymolwU//mSXZ2cCMaYYFYlsr0o/3HnnwVi4GGMP5LJg5GD5gFJBIxuUVLJ8yS+7iujg+DlsCAWeuOXNYASnP+kAEIyvNgKTU5Ng8ZpGirbzUmaRvzyN4r5H/B5GmCCf/yQir8djBliFISq7W6wWCD7h7hyDhrjPVGTyTqc0Q0YVYFqVXsPQhaAkJBp5CD5gAA/QNJAjGxKEimQhAE2hQbkLecfBrAbRp5BjgXY7CD7+QhnzBeUcfxDA+bTVoVekTPqtXBzDGjfBLjAC0rcJS+5+EgT8IKfKpAOK+Eyhi9qFw4nSAwhq4jiP2yAkZDZYQ0LGMUoxjCG2+HkHyH7By42Mg4IHIQOUlTJLcCADIHgagTlyMs/gkBHkDwDHSj8xzJw2Ec/jsQBf6QJPB4nSPXRhAsHmYU2EmkIQ+QCGEH/UBJGeFC/fxgjS0LMhSGwkqIRPEMXdkhDTchIRl3AASc4YcVHQvYnmvgiHAj7xxXqdhA+YMWR/0jBCEOYAj68YRe0aIDNrBcaVRxEca9JpCIF2cyQnMaZNoFmhawRkkPWxA/tO4iBtjGLWYxrI0NAxkGoJqR85asTdFmIcMbAA5uQ0YojISMYaWKHBgIQDBs8yAzm+I8MpOAjnPxHOVAAhzXoESFeyQkkZrPM7UXTmTZTE0RVEguKbmSZCOECF/yAG92MgEZ8e1pIqNAJ9XRSCyowBu1waANJJOlrCBlCxD4ShBHs4AGBUMXGDkIyc10UQ3P4CPqAOhOPFHUj09QJ/+JcUq0KTUAO1dLNDIJAozqCxG4Qy4ABOJkZ3QBQJ6ucjVhJJQ4l0UimIsnVA3aAgjwiFKkT2sA/UhbXnWQuNSr84yhbOAFe9MBQVA1hSJpwHiWlAKAGE+gIjCHLdyIEnq9xJxlINUn5kCQInCwHWQo6zGJsBSFWOMgx7BqbGDqzAOYzXc4awFeERCIoE4XN5EBCgDtcJy2WCMJuERIESYjnH2QwFamKlLYmkKEKWAkGu8Cas2+EzAymksRuJZkFXoIknQopRxRqcVClIgQIpP2Ha0tbXpnkSXM+FZ9ri1mZmcj2NfD9R+cQYlvkGYJvByGeJK8K0INk4aX/GIM7bv/hDvc84xkLQKVLxMggcITgaUOIZB23qhJOimUHgUhFA06jhdX+Y1r/cGVJUvEPC5h3JAcoailypig1gHZNA8DARm64kfbahAkyIapN6HsQQtxWDSzoxHQMcNXeHsQAaA3hEd4Cjhg0sIEhIyvIIDuht5yHRhWm43UxgtbHjCXDcaiFBUQbkhFjixs6q6sfn5CIkAQSxXG2yQTC4IlP1QUYlh2sSGgkCcoeBBxinHLOtrAYf9aSJpx8wKJHsAtfTEG0Zd7cgBKUINXEZCbea6FCkYkQOP+DxXIWdUmGVYcz6O9HXHYJDqr8Dx5EdnFKpklVB6MQhwTiSwptFE++BZv/7F0rWAfAhzNh8IVRHxsjJ3DJAM4QCDdMIRZDPoiRaQJB8QFUz9TmM7Ufo5wdsIAFS7CCaD1cElNwIk6cMIXhUFNXTctkzSSpMbZAIMgzI9slNLiDS+qQCkKMIBaWsJue9UsjKhAcJIKGdVy7OgU5ymAE4y43cWRzWnzr7MMXX3Y0lS2TODwjUkFQNUYmKeuNKIaJCBn0RetYUqz0KAcXWMIStCBpkXDAJu041oKioHEU95oncP3IvHOmV5EQfSOfBg3OP6KEWFB1OiUdOB0jacdpb0SSH1k5y/MVBA/aegRMQI5CpyUhkDD9H2zwOUWTKZNTlKTea0eIAIpQhK3w//EnOksDCqIt8n+EygDgpIK2EZLkfE2njiNXCS7EyPjyRf05PUrLuK2ghkmMpFjZ29wTDnJUue+RJtSIE85Uo3Se4H1aeIUxSRA3w5FoINQ6eehB0kCDWFCCCgboRJYMcFZZ11HbRia8nC3hwUU/gA9MEHcOLh9X/HzeJab/BwIYypGQWIAzFwENE9QkXwpltCbKAMLqQ1IUmcS+hjV5KAMIkYZLRAH3vBCoJcBZeKtvWeR+L7Ids64Tera6wawtaK5ONqru5aagBPhgCXIAAATA7D5i9jbiEOhKZfZgQlRsJpwlTo6h7YLCqVQjxw6i51Bjx0ji3mSC4kAMNCwONv8ogRcsgZ/+oRPqDyPspvfyDAcPLs/kRm4OThKOQDXsABu6QWX0QiEQcAYYMADiQHCA7SDAD/pcAqHQC0Muz9iiECEsLSgsQHGIYytCrHxiQUnwQg3wKwUsS0mmAwcpwB22oA3dIRPcYQUowBVc4QZcAQds4ImCwp1CAg0BJY58pASqYQkPak7k4B8GYHOQLlqEjiS0T+Oej0FcQQuDgjgozgKusHyiwA1iYQmyhA8ETr/sL4SAAQPIaBqmoR6aoRlAQhiqKCj6wQxcYQVqsRbr0AxwAAfMCkPy6yAs4eX+QQUc0BAbQBCIYAAGAAqxsCTgyg+Q6j+OzfOMzpl2wRP/gMgKfiQFaHDPek8chOAU7OEfzoFBakAk9EAPBkEczik1EE8krqqOgmEHdmAKAqERNmaYrkURlYUN1A5bMFDjLmAjMkMTkU0LKO5OEMLzyocGUAAFAsESSmAEFMVv1JAUe08SNMEfQEIP4oQezIAX+cTIKOGm6rEYDPEY/SBP9rEm6orzcsIFoiXeyiv2jo0DcC4Ca2Ihuec16s0CcuECIg5MeKH+RmiDgIECWDFnWO2y4uS6ciXDfMGgjnEftUkmhk0DAFIJamKu/FEK1k5RdkK8mPEgNM8lkIM3Tmw4VIKPbI5PQIAqYhDqsKr3mmAdVIYeDsLk4uSsZPBudiAK/3whDAigAzqAJQ/iK1XCBzAwtWYiJucqJhFx1CBRJaQPIcAwKARSNnIsVNaE3WiPQR6Aj7TAI9AhJAoJNiwgw4QIt1zQv9YRIcRBHMiAHtCxT/SAHCkHHrljHqPgFxChFhBBOL3hH6qJQuaKLOPkJZsJHkoC7f7hAyjEITIuTgLh9oDjF3cpaPwMB8JBcxSPQhAuGNSgKxKBF/zAD5LxICLgIz6NBWHyICBT1CCRMklCFmADRHbCH0tiOS+uIMtoNlYEBKIgEfhJUShBOzFipP5hEyiJJgQoJ5BgI9wBFqMlDTeCD2ZgB+ToPJ/RKjHCeA5CxX5HkL6BGbfC9Q4iBP9Lgg2ecyZILygsEzUKQDND44UqJBcyVFGC4QhIACR+IQYggT2DZSO/8yM64ZYmwQtGoANaYAII4SCiwa5caz/lDgiQBiFS9A0iBxOeoMdcVCResj+bCUZ3YhwAEjZA4MTMYgQQ7iOGNFju0o+iA3n+gQV44QNK7B++a9RutLSg4R+ECiNqNEsxQi1To0x3As4qcSRO8CA0swcmECNKIFJ4wk93Yliq1FBXJBD+jD1tJyTg9CBiIE4e4R804QcEiS8WohoCQQdE7JiATpAe8MZCg4U0TlOjJSVIAjOLoSTypDZqwnIyBCHCsn3AVCRIdSOU9SB+gFkRog//4e3iJFr/F2f4gkFDy6EaVKAHfuEa1PSi8Eo1OKMacAgVQmIPCDU5Q+IDN+IBMeIaCOQzd2JIi3Q9/6EC1nXPPkJrPGizqiEKemAeNU7F0HQk6nRzYhIkVrSZruk1qHAjUEAlLEdKMeI9VaL7JupDXWIBRFUk7PUghKFPEhOH1ANX9IJHlOMJWGAZ+1QlIkdf8a0BgOJdRUIDhmEn1GRj46xaQeO6/IsnaAQ8+vXrFGIGNgBn/0HnRM1gR6IDKUeHYjY0DuozfCIk3sEVmjPULlZq23FfbQJoa6owTHYtjtANOGEY5sEHZvIghKhrZwIzSUJxnrZC5tUmOANT+sgNPiINyMua/0ANWywI2UYuREviPApXbAdvaJFoClQgFkJhGDQgZQz2Ap7A/BxxNt7NvJaRbmdCM3HmBQ4VJNCNJ3ZAVhFiZ3ciFspVNqw2JCTzILi2MzYiBBk2KNjTYwnkWc2rqnoXPKiAk3JjBrggbX3gPXPBch3xG1DJUVvyIM4UIzQQxcCvc10iB0pAthJVNizgdBFiWGAgKPZtcWoSI8irM2ciIf8BNkmWVHHXGSLAGTCkD3fXfA6XJHJv8PI3s7AiLaBhHqAghk5rAioheYUOEijgBtT3NWS3tNKv0/6hel2C9O4kfTPzI4zNdD/iGVXjDmAWNuKgEVxix7iWcGjiDiqYJP/e1xnoNzaetWcF0NWcCX979zBcDjcoYRU0QHKz0gQGoBJyAQWGSXCA4h6EgBBigQs4IVcrBDkpyoNDgwnUNTXcViaicSSaU1kAwXUnpHt1QnAZJD42Yrgw4hPA4BPiJLFKIgtIIsnaOH+BIXhngBfiYRiMFx9MYAL2IBdAYGOAokx+IRAIYQZmIBe2YYnlDAA0MW5tAhNSMLZkYzkhxHaBaosJRHtlIn5ZODbG6R9IwQgQwgjO+CBIASREmULCdiNoyp9IYoNESOTwFxgsoRXwIhdAQW0ldw78gClAAHDWIA6E4BlyAThm4Pb80SwFyYpJovkWOSeeWCfw7m1VopL/S8L0WpZAcpdBSPkjzlibEeITuplBAAqVZyIDaMpWgEGEiqyN0fkuZkAb1FYUfGAOWqASEiEWzoAcCMEYYmGYB7kVeIENlLiokjkknJmZacKZozlnUPMgoCWhKwR+K8SUEYIdSKGiy0eVP+Jwz2OXdimdW1n3hpIoiZISKKEVWmEGysAqBnmln848uYADNsBuYyMzyE+hS0t6owXTEGIo5hbZQuCTFeETTOUenGGMDwIMiBBb1vgjaCoLaOqfOjqdRSgFLCFXLAEp9gmlwQSlMzRDDYEPwpoXqJhPeuymb7o+bUJQ/8GmbeILCPofgucgkKDjKoSMHgEX7gFKDuIT/0JgThrAGWxAlP8ADBQBgN7hHWIYQ85DlTNaHv5hjZ86qm1lqm1FlkegEyhhkFX6pLt6BoLBEFIgA+6DD3ghVxLpkGOjraNZTUX3rPlEhybADUAAE3bgDUCgCMB1JEjWJhLbJUz1Eb6hGxThHwg7BLDhHx5BuRugGwTok/8gBrDBt3einDNaJJh6I7A7nA7inyZbqreRRoKhFbz6sz+7FehvH6rbEkqbD8Bi3V77Lf8h7kiCBbqYQRx2cUJ4NnZItovgC97gC0DgtncgFi4gF55GQhFTJ0wVF6a7JN4Br78hBIibsLvBRBMbwh8hsG0BrBYuKMo5JCLGqVXiRoZAsv9TYAgQi7K3EQZnoBWQohNmkBfK+amfWh6YxxIsaiNOwh9JF75nQ1xjw7Uppwfc7DVQgaFnYky3aQL6+7/fOrcJ/Ak0s0IbiLdlAhv8ocEX7x+QO7nltBu6ARu8HCNwQbmRG2RR47FHAgizeyTWfKbKWbQRC6DG5WhaYR8QQh6yYM9r/KmJRMcxYqZ//DWaDyEy5z//4TMHnSSkWFEpZxLGEiRCoSTgeiQmgH0+4Av+GwAA/A2UAQamnPPUCCHqekJM9R9MdIz+wcFZndXhScsxpM0/Ys03Yta5Owvi/CA4GslIJzoyoM/5PAsK4Z94YQRuNSSQdTaO2efSuiR83Cb/ajQzTmzIVQK/W4jSD0IBkhwjLpmZOOofDsECErnT8eANdiDUL6ASKEEb5lp80jy5GUS7gfDWVeIIgDAL8j0Dcp27ESIF0gnP+WHP9/wIhn0buMAjkB0hMg/aGYQD1C21L+6gRzcnOK8/1bLaAQkjHBhbqHEjsv0fQH4n2k4ZQCCR8WAX/lsZSiCKnyC1fifBv/KL+ySxySjWDwLV+0QMaILe9X2N/0mXgj6E2MIS5EEetoHP+YEfLIozFP5AOIHZCb1Coj4kXvICGhMhLCDjSUJGlWW1Jz3kVcLARUIyjXzuJgLAWYAPnuAJKiEF6CAevBMh4rd8UF2Tg4LeQ6IN/0Ri5zFinO694PM91zPAfv0pA6zaEHhB6fkhF75kMzYiUhhgERYB6k3BQD5gCjLj8QmE6oXcxHRmWkIMtlLDohpzySlEdJ09NJRhK4aVJM4gJFyvciURI3RIEXuACPbhBafCGA6BErhgCLZBG/iBBPLgHyS0AhqI7jcCm8sr722Ckw8i7+/d52cKsuc8C6r6kYiyBFSg05seM3bgDriAATiBA0xhESyfAz7Acc3TEiydolDY24Eq0AHlCertIiyCdVMjmQACyL9l/woaPIiwoICEB58wNMigYKIeKrhkyZBBXpZtWTRu+1coy0OGMUY+xGUyZUKUKlumPHIQpkuGyP8QHrkZ8mKWIRh3XjySwUCnXLl4Jcr1b8SUKTt29OAyi8OsfxzYsNnHixcfoiN2zPz6bxHYsQ9f/DNrUAKffzLIun3LMCLcuWC90m2pxW2AfwH2HmSCUEVCLhMKvvjyJtcVedsyXJSH8OPdhNj+lfxXeeYjgywnf5Vpsg3CmqQPthFT8+aRLDodu2YtRl4GXpY6DbVUlBcX3Vx2i7OUdQilXLF49TD4xXPBwsqbfy3wD7pLBHS5FBTrPLv2hxbGhjobKUB4vwjb/oPBEMGAf0SifAEBwIK4VawzFIS5rTGvK01axlhw2UzEbEegc2IYdBNrCrKm0U1iPAhZBkPwkoL/JQbwYoCFKcgjDzPyDEEUL8YAUKByb5SYEnooGkTdii6+iJAcOkRC43gBFPFPLCUUdME/LBTEBQPU9bbeIS9g8gUAbwAQCC+rQGaQGLwYgkYh/7jzzwIqRfBPBM7A6FlNk4n5j2gjmXmQSAWJlIVqMInRBj/IwPkgP3HGyc8ReTLDSy6J+KGCVyCASWihcMn1D3VuGMpoSwSpJAcKNYrX1xcSwFACEzI88QQLFhQQZKjqcdHeF7uYKgAAAgRiSX7IgBiLIZ0MAQpYXjbqlhljukXmP/JYqdE/oB1YJjJtGGsnsnEiIw9t2+RiF4HM4UrtWAMQJtd61X5FnnMS/JPD/0yRNkIujeJZWkIJMmzKhKcFXBsqF9ce4t4beKiaqgp80JZLK63wYUkGoCHE5bbaHUhsQgmj+VWv/4iZ52ojGYsMBKRBgHHFxoqRBS/MbMNFLHdhktK00xqMciPpnYxytQKl5AIR/5DbSI2RvKHCCCzo+IQbLBRBSG9CMzABqT2girMbifDSSix8tDJDK5Yc5DBCX5I1RsuMkvlmQjAhgwwJoNBBAgkQPIzxw1dsw882Lf4Dwi5xz5XciQ+xXKhgBK6nLV0yLzcTerGYh5DdWsNYbo145CxBcbMYFcshQzAQLxfbTHhIVn3yMQMfns8QjCEpuCRFl4efnlBNZjKMEP+xCUMAytixQ0DCKquweNBCyZGFlEl4oz4TAR+81W1zgyIk8kHH0yWCSQu5GG5CnBi0iAcJ1VxzJF8AkYMKLPDyeFYt8IJV+VlRkkgnlOzRib/+et7K6AdxOHB2V7cUwWUFF7Q/mA6fDRYAKmxi/wAgCf5RttiBYhVz4ATIQhaIphgOD9JiSBcKckHgRWcufomEBj9YkBH8IznDQwgCsHM9cgkACCrIWQ9asJvz8YISM5yhJSiBQ0q0on2G4IMhKCE/+4AwOzZoGZweIkAEYgxjV4AAP9o2oQntxgLPK4hD7tI3upBIOTsai3RGCJZueVA7hCuI4VrWHbr8KD2JSkn/IwSACQvkzHu80EZWMsAP2WAIOJboYx/vmJGNFESIkIESgfqnEmcEKDshaF6JDojEmZjJbJRcIgSusIoMiCM3hzhjSkxAFj+cTgWeVMnfCpLFhwDCIMVDCBwKgoKC9MAYKbHbFhmyPIOxAAbHgZtBUmkSFUmABd+CCyZ2oIwW9iAQseDCbMSUtlXw4x/TlBM1oaQml2RtiB+EpEGqVhA0pc0gZlsF7TDGjwwAZwhcCMQbklNFQ81BJXgAQfJMEsuRqIguscxnoShIolImJJfcZIiKflRMsqxyhEVQgRwdugNx5KeAqQObaBJWP5Vss6AcfdiZMFbJcmIsBcAQxxAC/7GLXfyDgtXihUoIyhB/FuiUCaFpt1r5lVuy9CF3mIxkEuICuCQULL44SC8LkkayBEAAX8BEEVhoARAIwAJV0AYyzFkQb3q0TAVdZEffwrCzifWcId1GCnRjjECAoJTxbI4c7rI7k7xBpf+QKV0I8NaCEEI7cVDJLnb60oPYlT0JOSrKLvGPthoELSrpq0mKYAELvEEAIMiFHMQRijnUqiAALE1GX1IQdhAqCV9NiVZTAoE2jBWkZEUGyDgxAHEQQRyTqaJit+OJvJqEBtkhQEFK6BzHMpYhAigqXfEpWMCOJAooe15R/yFQhHgAB2R5z0oDAAJCEIEA4hCHNuZAh/+zVQyAbcioIa3kK4NIhg6lpctpb7cisY43pFdwLSdcStvczWUhtzXJd+ByHN3GNDs05etKwfgQARz3IYZlKQpY+gyTGNYkAi7QcwPw3Ak/BJgpwcSJFiJTvOIVB5kFBXkLIqYDWUkkkqHuP5xABhyQgQyO1KCumkMCssHIkjy2GCgaKIcCF0S5Sk2sWxIwlnhWeCSI7ehwEUJkgxxHw1/R21g8AZZY8tYkx8OwggernZ36VmZEqEId8KAEQgzhCiRwWCGO8JEZNyEEmxCGFKTQjHMUhLTVqsFDrPePbDYMibTLMR1AccArGAS+BzmtSbQqVrMtEWxguwIdtuEJ5v7/Y8l3ea5BFhyjr4A6Oz29Q1Lb+xBNn46lo2aIpwlVQt/+gxBRQEEsdxGAXURBHAioLzWv4IpMNONL9yvIOfRsMD8/5KdtaIOaZPLZ0ojVIEksiOxWwd6DbNYltSrbPxBdtkpeEqSr2MYzBBAeVbcM0AkJxIqo3F48BIKxT34IcPf6D3e7Bcst8WctyPKGQJzhRR8oIQWG/I9aFLWo+XyBEpRwA1cI4x/F/geyU7JRFCmbIewuiBhmt1WDmKk0qh1v2qqtaAjQYRVVeMY2sB27VdSudghxtLXDTQI20w4ZC9xGFXBdPFmjmiythksJgVsocqXkBfo+SJMRgnShf+Xg/3D5d0twOpK3eQbpCPn30/GQTxy4Agmlu7ixC7KCf7iCQLCgC2RkAoFVXBUUYFMJj3POWnIWkA5zGEIVxEGBIWzjClfIAyjyMM+C3K7bhjc8HfLwijzwvdziIEQgttiXvZDHt1I3SJSHbhIlDNQlGDgIFrBAqDjEwRoGKYZBEDvY5255O6X/x9O383mTdH4yl3iu1REy8H/ggAJIYAg90r4iPejBIM2oQBL4PJJB9OMKw3oYMvJwBU6sIg9YTaJowkrW8Idb5ge89N+rQAEKEAALIJB3IMjxDAKQYRUJSMD2RSACwlvpGWp191qxDnrKUW8zgXqlh3oBOBlId3suAv9mnlEHBREGB/gPSvBviJASN3ADYrcOzvADBnF8LtIMKdF2g8AQIrANbnIgyAATYrMNDqQAc8B91MZVBUQ7SkRJOIdzq4Boktc8lddygYBhfrELVWAQLlYQ1HAQyZEcO+VBY9QyEjgWiLWAKVGB2YFlD/gQUDgXKlMQ12AQcbBQBvF7olcQA4dYFpgSWjgWYWAwN/APbjgZWFgQEYaGCRF8BfFWrmAGEmcQE7cCNVAD9EAPekCCCFGIKdEN9FABzdCB/9CIMxGC/7BxBiECHiB3IXETeSIsJDAHV0AGCIADhfBy2ydzCZFyNzhzYqODqrhAC0QHCTAEA9dWB6h1CIj/hHDxaoSCBWzIELtnKAN3h3WIEGrYHGFYKGv3FugAFy+Ab294A2lXAVIQjdPYDHqwAuGQCSuQdoeoEpFIF1cjDH42CNRADYGAAmdwAy9XX0dgUf+AfduAAzggeOKAAShADk0weAvkTWeDijLnj7HzeHRwaNrgAfmFgCkhh4XSgC2BhQn5EFQHF1w4MwmRBv8ACBJpEjsljAYhh7z4D0XnEr+nQar3EH2FDr8wFjpgEM24dq5QAQXxJdFYA66wAi+pZ+dQAXoAiCPIZy/piDDpjXQRgo04k/+gCRz5D3+HA7YDCph0BYzgBDggDmRAj5dglbimYOTwd2s2ivl3O9tA/wZDQAHiUAUEgH5Y8AGoF3yeRgMeeZD/IAioRg5lOERWWRAbWRAOqZIL2RKuNxOO5Rm+CBcWOHsqsZAUYAaZ8A95VgErMAjQZ3EGcZM+aTUE4gwV4AyOSYK85U9Y8AxhUHpk4ASDF48YKA5Y4Au+EITFoHAKh2G2BpvmiAKXUAsBoASg+Qyn9w9seIcGkYsuMYUqIZIzAYcMMZwMEZdF5psa5JCGYleqsB3NWSA0QAMqCUuFSRYqg5EmYZ0HcZwJ4YZ6QA+u4GfeWHEwCSaU+Q+ZoJg6sBfB55GCWRA0UAusGQD1iZ/F0Hs6gAL8CZv3+W/J+SISKZ3/4JcTCRcAWP8Q3QkWv/edbsGgLSEEb/kiF1kQq2SM/wCYI+ENBUELBnECB4Gdk1GRCYGGNPChCPGbaPcPK+AKeqiY5imZI6Ge9vMQwrACgtChCFEHbnkQB1d7e8GaB2p71WkQ/ml7E/gPBZpwKNKb/5CiK8KXM0GkLzKhL/JKZFGYIeoSAtoc2mmhFgkIgLChLZENtJANB3ECKDmf22ENkACd/8ClBxGnsFRX9lgQGOAKYkcPi8l8FBeZCVGj5wmoI2F2X6GYaIcBdUiGI4F83smaKkoDKFCYI1oQoiegxZAN2fCgKmGpbWoSKnOmaVoi/fEV/+Z61lAMVdoScHoQEWoSyDgWcYn/SC3RAA2wBgxRoi3xqVEIJloyEsc5pw/xqC/SnYKAATZADRI3cQZBqGNROgcRlDX6pyEYrQnhh/9QAZlAAbwlBEd5F663ol/xoaz6EBGKCKw3E7D6ELVnKK5XC1bXqS5RmIPlrm8hCEoArmOBq2uQpQUBB6/UABR6rsbpof/Wq25Rkbs6E9BJC6xZCzRwCSdQOjiwAke5fP+wDspBrX/6FT75kn5GWhUwnjpQhxN6pYXyb/N6EFsAohD6D+pqEo8KkS6irqogkazHW406FwnLENfKEPtKFrdKF5AAF1u6LThLC41QpwyRqIVCC7XwCzQQDhY7cX26sek5FhXQmCuw/7Eb6wpbgAiw6rKTWBDuEJfokKG1QAteqBIpyxBR2hIWWIcW6LYuwa5aYw2qkKajGqdw6xJzWpikmhK1CrgEMrBjYbQMkQopAZ1NiyKn8A+QALTNcbdfwbAHEQfcYBCqsLfXEAJmEA579g+bkBBZqx0X9yWH2rEGsQ7C4ArdYBCNKaf/ALguixBPe6EIoZ2g2hLFZxAZqhJ4Kbczoa6rtJ0usbcYWrxuwaUqAwjocA2kKrwMoYwmYYG/MKzDyz94iTqNmxIhur0wIg0lgghuW6YPkasuEQfogA6NNBKo27pbOxIZOxOUuQ7dMAjCsA79u61iV7ljIbNQSrdsyhDA2v8SuksgYTjAYJENqnC5yqGM6NDAX8G5UMoQ3jsSPPAPp/ADi9syujASrEAwjHu9vwDCBXG4BgO8zvGvBsEKcJAGcGAHcDAK7OAEimADSSCyJjG/nvG1H7sOSdANr6ux/5AEyCe0B1F8pjsSEAy5kAsJ4DsSBuwiIWqBnOtYjtW8KnG96NDFdBHBbjHGXBLGCQG+i3sK0RqCtYoQ61si0dBXfUXF/9AZDxEBkHsQAcw/D3G3mZsSqeDBkmsZkxGljgXIKvHCdrAGJSFa/6AIsiq7ztGsDIG6M2G/G1sB/HsQpCUMbVd6CgwXdYw/dBGnpGwSKfyF/+CFqwSdLewZAez/xCNxwaxcEKqgygmRvrbsFgjMEIyoNdJAxTFsByYhuahcED+cEKs0xi3BsB/MwaTzl2TxSv9qByHADn9QEH9QROvpEvbrFpdMF/1byQiRBDQ5k7j7FlQMnaicCnpMF8iMuQcBDqxcvXABCYi0wndJFlwaAeObyBIKiacTDQA7EoPcwT/AA4RcEAz9EJJLyI/oFi9cECQMJolrEg3gDE5gA7awzYpgBisAmQyxCWnXzRw7GeVMxGo3COy5ng7tFiI8FvLcEqzQuKlg0SqRywhB0yZRzzqtElKw0wkh0w8BueX7D7pQy/8QzSqhzB+EC9FQzAeR0y7BJQUDwj2dCgHt/xJIHQdFvc4uAcfq2wDhAAYH8Qd/4ATIZ7YIEQ7JQAot0b8MUcnl3Id3PRabgLpnDZWu8HyZEA5p58Z8PBNpUNWp4A8FQcW7/BVVPRblC9YzQcq6EM0/ENEuIdH/IA2swNUHMdQVXaI9jRClg2eEzRAokdOdjSK5CgdrMA0P0biODdQgfMeKbdiqrRIFjdtj4VgBOxO5ygMgbRC2YAs2ENIusQKPbBC9AAYeTboFsbETx2eom7Wk5ckGMdLYSg81cN0FYbqbgM3/ENe9kAzUINLc/Q8uK9ER4MYmQcKoXdEifAqJ/Q+p0IE8INvaQcKsgBK4kN8aOhb1XNSQ4MEtgbhnBRGUBREHnN0SDI3MFG3TFd0Smf0QBX0604DR/zDVKVHbCXEKHW4QSJ0QrzTWI1HQurDbKUHhQzsGTuDc/xACxZ2Y2T0Ssju6I8EOcY3ErovXGpsE62C63f0Pdn3X3bCHPI7EilAQvVAQySAC/eAK9JAJ202TRgvTjZUQNawLcMAKrEDI793BV04gcBDV/wAH0lDNZo4Q/03UFbnUYJHZ0oALFL3KDx3bjm3hBSHCJFzQeW4SMRAQACH5BAUKAP8ALAAAAAD0ARkBQAj/AP8JHEiwoMGDCBMqFGhn4b2FCGsVFDBwGsSLGDNq3IgxgMZQiwYe4njwG8mDmHIgfLEwwUmBJf7FFPgFohyBN19mnHASiM6fQINqDDlAqNGgFI8qVXptqVOE3mpFOlnToKOnWLP+m8DhHwOtRteAHfuvwUI4ZNOqXas22z8UYwT26KFihAoLO3ZU27tDmYUpgSwEenHmH7lD2zgpmHOwCAuyFi+iZQsRAeXLmDNrNWu24DELCcVWVXhHbee1uQpWG1hO4KSEr2Mr9VJuSqwnJVT+60CwaFAZ/8poHg72EfGLLoCKDQpIIOfj0NN6+RlAAABlYKcXbC2wmoVcXKKL/x+v9gD5i9wIemyutelUguzPDxS7PHNtFSoQHis3qRoAgf/9c0xQXjywjEAGlrMMdwMpQxtBKnDBCSfyVWjhhVrVh+FxEmQkwBuxsMCgQCMmlMsIrBFUIkLaQYTdP+Uo84BAMv7zQDkz5jjQjN0RtIsAAkQi5D+eIBDShiSFZ5QoAmkQVHJIbmTSQPlFCRZvVo5hTCAatTbDP7FMsd1GmPBIIkcPKMOdmASx+Y+bOzr4T38C7fBMRsANxISVfPbpZ0YBQmRcUgNq9pxaUyyBoo0GvfiPozRut8NAauCoIolwljNCMP9waohAapyp6T+GjACnQWYKtIsvf7YKUQGuEv+0RKzydSGQrRA1QEMPBVxQyUAT+BFsC/8QocMzLKighho5oBjqQlNMAWlBD0xRbWvVjoBGMMFoawgVaAAjiSTd6pgtqcEEwmkVA1FhwBC3UCEJGv+AOxAaQxTyj76xjKBjtAKJ6agyPTAIQCCBjPHLaZk90oCGC7Fhyj8cfHWcS7RmrDFHhQkE3Cz/JDLCov+EqpLJ/6jAAh8EqVGlQVPwQXK2VdxiMxXcokHFP0NI0sQ/ffwTwtB9NPHMFKMSBK4kKQxRs9BC9xHCLeNS0YS7ijQxdQhRj/vPplQMAQwVMyyqRi58TDHCzp3eQg44DTz0EMQXTkwhJ4REZ0LG8Az/d6CFHhX0mEIPCQTDZRPs80QslLw5MrwC9XHLop92W5AKahvThztm9ILRO+/gAocuMZBDjju+xLAA0CGMsgAPuvzDw0JDIATGAjE0IYkiZDBSiAH/BNEJp+1mYEAwX6JoTDDPNBGDQIWTxMY/FK5l8cbYZ6+QR0lplKdSpRXEBQcgCzQLF/2SfFATP/9RCDACAQN/pyWnrEIV5FwUO2W6dGOG7mSoXfCCQAVgZCAD/xhbEILwNTFtSRcN6EwxiqCRrhyJLRMTiJK0h5lSCMSDHAwhQjY4EGbwogRW6BTwDjI/g2QhA4Xog+qGFgJ39GEMGFDCP2LHCoXMjiM95IgN/3zHM2AYIAXyWKFCDKEGMY3gGQtrADpAk0IRWhEoDiDIOE6ShisaJHD/8IlAxLiQPWVkbz/pCgeIQAAWzIASSrxICw2yv38EcYfQYeBLgtAKU6lhBMZAwWNmpZvs/eplfCKjF3WCyIyBECgUQgAhFlAFQxgiBZYIxiUFUoUqWMIAc/wH8PTIQisusGxTKAElLhCTWT0LHRuhAR7E0wOZRCkOA+keWLIonihEqUP/oGBaxIKWWGgERLno15c+mQKeDUSAAwGlDTCgCSlUoALCEAZBMFCDFZBhKTZwxTcFQgYjUsYSaDBVKp+QA0z8A5aLNAjD1sINbyglULoEi93Icv847LUDKxZQwSH48KUZtMIA70pICsRBASSsYy16KAg9amAGcSBULUqMY7d2AJhAoGMyBbFMPBOCxn/gYKQLoVAGTTE9jezBii0iC5SI9A+6/MMYvJjBTC7ZtIQ8D6Ua0SMDcTaCctQmNVwg1kB+UdN/hOIfIhhIHoBKVY3tQiAg+EcqnvKay7DkH74USFx+4g/jVBUj9EIDGoKwrZGpLRCG4EI6hvEPuvKplkGZ1KSyF1YLlfSs5PkpeZpJEMIeZWdUIOACEYrQFBigEzMoWysowYyQAVYzihzLBjDyhKf8VSgXiOfq2CLYfzjjIN1QCzQPuJAsFFYg0GyXQAywM8b/DqFpKcjAEIxniBkQVBzk0MUaplSWBtijARGQgws4MdN/TE8VazgNSAXyqz6NZiDuDEqHvrqRZTxAC1bC1WWRZIt/dGNo/yDFJ4wgEEXQ8BPr/ccn1FterlmpmcCrXTNve9sDHvCFGbDEP/jAB0rsgxfioIQlLMGLf+QisjNAHkEJWoJcGGMgoMkKNNKyVwDM8h+YaOR4yZJVp/DITO/Z0GkJEgGjPMIf7/jGApxgBDD8gx0hMOs7BvIIbOBiINg4SiFcuxb+puCFSM7CNv5xhABrshX7YAYzMiCPDGwjC1WeMjB4oY1ZEEEh1W2cVnyglDdk+DxdDe+txDOtgihg/yxXDdQ/LgAriLQYM/4QyI+DrBR57Isgfv4HP5g8EDEYxNCHNsgRDkLk2mXghVc+whHEMGlJyyMFneiEIXKRAlCsYhvbYMOEONDSUwmkkZSABpMQsleFSGzEJLng9UYMTFMjpLlHeQMevvAhFcSCCU94AhdMIAoHHCCq/4iLEC50Z9NmrBCBRsY/2iCGNiCjDfygNjLEwI99pIAKVOhELjpBCXFvetPkVjAlKNGKTkw2PI+EtbyHM7ijdJYgCGCASAfS1130QBzi+Ecr+DDwVrRiW4bggyGGwIjUIkEgD593WqTdhn+AAhRXGIi0BdIGCHQcGRC4drb5gYwjXHsVvP8ghBtSU92sIMADY6k3ccDYKixhZnB4PYg5LliQ+LxJAh1iQSzu0oMBDIALR0+6H3rwAhCAYBc/AsAOcsELXhBY4Qa/JALlkXGBbAIoERjtP8Qu8YuQoCDI4EIG9tF1ZhAAYW94w1V38YabGvPeB3GJJ8hT94Fwt+wXqXOF+inil1TpquKQgx/kwIVV8APBKVjFP1YBAY9DQAyIlseiC+JaIu9rHsnG0BgivpBlC+TsG1cIBE4PCjrkYyOgMHtCVl+Qs5Pg9iSAQO4rn/tVDEEcsxDHpGJxm4t8+B/XRekNNHMJufyjNHg9Pkn2rRFaCAQQbvmH9F/S/LTQfCBfxur/P2gQCHFsIw+x/0fXTZoJJDTjHP+Av2nP0QyIex0zsCDIIAjiiitsY/MCsXkACHKggAwZ53EXsXq6h3tnJxBT5YB0AAV08Ap0EA8P6ICnd4EXyAi19w+5l3v/oHsQwAi4BwokcHF5gADkMEvNN0t4sAvJ9w9vhmw4cRDbhz0U8A8f8A95sxTEhRCX0ByN8A8pJhASgSGXkE+ucgISEQCsYhA4cFIDcVrw100EQQ39IBT5BwvdRA/xVwEFoQcTlX8IMQjU4ARXsHHSVnL/cG1u2AYdV3HIcHtV4AuBUAWFsAp5cHa014D/cIEEsYcmuIeESALoR4itlwzx8GYCQQ3//+CI26MeAkEIO0gAgHcZ0YAVOrSJA4EI1gcJ/2B9WWEN1mcN13ceXWQQkTCEBqFDCSGK/6ADA+GKBEEBEfUPzaAHK+AKmQCGAwF/8pcE65AE3ZQEwlABetAMYOiLv3haK4YQz0h/ArGM07iLK0ABStB8shgGWPAPYRAGN3ADhQBzjHCIeZAHekgCjKCHIvBpFOALtXAJOoACSkCPcIEC//CE3ogFYTAQ/XgQOWgQZhCJl5gR/ygUgpArZTEQnQEH0pCKmYgWkfESzdaK7fEPgIBLceBz1fcPR6gRGKARqWgQspgRNCAQP0MNrlAD2EQQzFgQzPhQCwF/UlAQNakQNf95kwVxDkkQDv+AjMJAAZmACASRkCdRDAaBjyU5EN1XEHVAi2thlEIhEUiZfQhBdmMBiwJBlDqRkyegkxxBN0uhCgTBVBujCuhglksBB2ghDRcRROkRioAgBDawAgNRAwkhkyShTS45EA+lTdSYEcNol+sgDHp5jYigA0iwbKSnEyfAlVFClhixBSTxcI35D3apEHfWFNlnfbAYcSVpegORCndEECcgFP7wAxx0CgsRcS2mmgaBDqlwDWSZCumRBiPZKibxDVxjAwPxB2ZgBnZpl3hpEHjJlwahl2yhnF5YEOFQA0nwD1sQAc0GlhqhlmQBCVu1nQsBCT/AmgOBSxj/Ip7vhBD1t5UCkR4NYSHRcxTS9Q/TtRA9tJ4XcQqlORC6wJ3/kIk6gUtumZv3qRG6wJYaEQJOwDXlJRC2AJyu8A/F6aALsQJmkAz5kA+eQwqMQAoEwQ4rkE0JgZwfKhAgugJm+A/RORDCMKH/QKH/AAX5wA5mIAKDcKJAIQ099GMHsVUCEaAFQZ9K0ZZwYAcECp9C+hPiOTv+cAr2aZ4K4ZY7xJ/hyQpOShA/hBDR8AhdFA04ShA+ahBSUJFgIZYKIaZLMRVNgRDABHhv9maoIBIvoQWFlBCpaA9P0aaMkQCfhREx8T05cAx4oITH0RUGITf/oEMzQRCseIk8R5AI/zFPSEJG4eMnMRgUjMGIJOGoBAEH9kQQRZgRMicQ4AURjKER8WkQciYQP4gZgpoTAkGmBUkSWtmjVoKphEMep9GeBRF+WNE4LMAm1ZBmECEbshGsq/EPXGIQSzAraaGssGYcDzGRrxqtreIGFgCsGWGtCvEg/9Ai3IoRDFIOKpALI/EP41oQuIYR3yOtGKEAlnoenaoUrroR9UGr6mofAxJTBNFmTqEMq1Gsb+AGE/IP51p2Tak9/2QeGhOvV4QxGFFi/ZQRb8ACtaQmMKKv/3Ag5/I104GvBWGxGOEF2fUP/wEAAhB11gEkJYuyPwIkK1uyAxEALzAAnABzlvgU1P+XEVs0HjAncW1arwqxdxaSDVklJjOyIm3SGqGSSa32KGaSKlmBHa0RtW+SEC/yN4FiAeJwAzrqs5fFsAxLELh6EVtLHtGwqVQFis8SRhkRC8GANEbbERTBILaGEK3BUQmBLdbSIAfhBf3KEWVgRlx7EidQroEbTxjztY06ECcpEGaUCIT7DyGJEGnbsYwCBNIiLQfxrTuiNuk0EF8iEBbGGjmCNEIXCNWgNpz0D2r1D40zBZpkKiOgcJawD2xzt9yxGpgQCHVEHzzAAw+xpRwxa2nRUlTVcuKxtIV7FHFRAjLQAjKjGyiCIlXCJjkQM8kCEZY7Ap8KI9ESC1XQBMb/oDafIhDgsjOK8A+SQAaFQDxIMwKfW7vkCww98w9/8AdUIwmqC27g0jM28w9UgzNvoikLNgKTOyO2sQOBoD48QK8bsqh/kgix8gV/ehQhW0cQcQj99FJZYbaTGh0kJDPU+w85MDhjNRAnIiYoLBCOMAXG8DTrhxHsIBC3MAa3kMCGwFbygr4/I8NAIxAhEA5NoAhgkHEcyAiM4Dn/4Dnh4Ax2MAbiIAlUkAGERQWl8jUzwECtYAgLxguBAA5rQKhmobAJkUHJ6yenKRzy9q61ajjWwwX7wAVUsCkzQAWWAAx1nC8CgQE/UwW5MFStWz9vYhu6u5488DwB+Q9LRhDO//BjPcQKuuDI/9AQdhBE9GnBF0EGXMMK/pBaAvEHQzAE4La6luAuUuwuR8QLFjYGX7yQUSKo/zAxwlvGWQGtQNVX0MEAXDALJ5JCIyBg9aIQkjAEtPXJ//Az84MwVXAn8qkROMoKzawTuiNABJRbhiVbpeJE5BAHnAFPG8FSHEFmRwG09XqoGBKnIsQyWeHKXcEAfsAHajADnRBHGCEvhdAE4PAP98xDdrSjPAoWOIoL9Bk2R5BEGZFYnVBUTRRIa4AOfzdGsuwqW5Sz9eoR2PE353EkhMDHxiBmwMBAwBNKsLYzljMCwVYCwrEEVZQ9xsQngPoUEn0QoEgZY4sQ6f9KHMIkHwTwC0ogDpdUKsFwURwxSvKsFMA7FiAtSgPRLWqzSory0D/xnxipFN+HEPE2EFcFFMR7EnQKESWmFeojEOZsFP+0FKaXC5SwKK1gCY6FEIZFAT/wDueZGStwA/hLGWyDBnbLB28ACGLs1OOFqRocitCBdxljDJYgMwLRCQ02ENWMvwwFomsxkA66fEetFNUcTQchPEFgKpOwA77UgyLU1whLFurDrHXzyheBznxicxrRIjeYFp8duk5gIT/2jMcRWwrRCm27rbURC89wNMdKEOCMJH2NEWe2MaFFEMdNHrw0Hl5wqovUYjENHZctENUtFGuVWEFgAGwlx7H/wAfMkA4C8dLkkWGpoT1AULBZsQFZrRC1JHgcdKbYaiGltRTPc98VYli4bRAI5EwYwVjvglsZgDMzQHwtQAkniath/A9JKhCnqRCR0aVk8U9j7ddH8Qr/gOHQMYTzfSG2/RSkYATstTGetxDAE+D95V+8ZVB8cAg6wJaq4A0QtAZrIAU3YQrakOP/sA+JwAcsUAUooI8aMdzjUXf/8doWfhHISx5Ljj0hEMMCYQS2zQOc/A8iDgaK4Axm9RP9/Q8ljhX6LeD+VQiPJsUGV2C8QAkzgAYGFWEsrsX7wG6pgTlpsWEb9qpdLRTbyxG4YividREAEHfEgbjRAaZOsWP//7DlAmEciJ4Q43QS+sIWriXFWTAEkPZnXv4PGcAL7tYJ2yAGkSZp20AHq8AJIeHKCBHYkORcAjtvAQAIpmgUNX0Rd7MUI/sPxaoUKpEjTgsWfvACFvAFb/AFXxDoJP0ElXABXFCB42AGWCkQHy5C8oBoOlFxGxHpiJwFktYGJncE2sYP2wAMudBu4pYLUaYN08MFuQAYHLUDZ3Zve0AJLSDe04ezSU5VoXoQyTGwRgECQCKyKlMCBOYHq5AOnwYMq+Cb/yCaB9FiLVbfl/HssUJxIQhyIBeCcdiG1oZtEEByYlBy/HAEIc8P8kC7+0AssxAPArFqZSeF53HVl3VBQv94EEInA0/QAxZgDFzABQjA8zs/AEv3dE/3BtaxA7GQCy1QdbzQArrNB7mABreQeqEHFKNl6OpKe7r3D3SAjrxXeRZPeaCwDcHwBsGNECwvECJwYeNx1SzRMR5z7xsB806x50HxBlGgeJywDVyg9HufAlWXCOU2boaQxe3GC/uA6dheIRJfECV8RWdHeatQ8gi2YFTHYIfABSOxg/LGqjy4EVPx+VkRCz2w0lYUqWqfFTkhBwSAANvgeJLXhgNhcgThWvJQCLZfCBnnBImcB7cgH5kgEKNgFFgPgqcnEBxocRJIB//AgVPV/E9hewz4gatAAvxQCFwgfILewQVRPQP/geRsEVb4aCXFnRB5nhaHPBDvgX3YU7MCsbjaNxDhLxD90FA/6WxSsGLNaRCN/xIPChD/BA6sMXAgLIMDXfW7UkjgkX9ijkhsI6YNsoFt6Gwk8a9NQpAh85AgCYqEyZF5BILamEccuUBkROShEy+eKDrzWtL5B6onyVUkSazKE6rQEC5ybvwjwDThroFQQ04N6SskEapZtW7l2hUkBoFhvFKVNtbsVKv/aAnUcXYqoalrrf2zNtdt1zP/QNzlOxDRCa04/uHA4aqCs3/CaqzIlESPnhrUBoXbOmjQP1iwVsCq8fhfM4HNzoEOeS6kHnqbL/+jZg6DEhS7zuC4kgeC/0CMFyG02Q3BN7JVEHxS2LXL1/Hi5LCIE+fhyqpVPenkeUXnlUronP7dUmI1QK20AvtNfWEQRV+BxRIGEove/fuEewPBh3+PvsAFZtv/qyMw/P2E1DurlmL++0eI89xKA6Q4EmrwH8CyWsvAf/b7xxXWXFmhgn9MG8s0D6cKkS8Ok3AliQpqoICGS87rb6umwPqHQF8K/MfAMf7J0SAaqMpLoLX6Ui+brc6wEMB/2hKLnLCQdHKs/JBcY6BoBIKjymnGguSfHiEM8pcnkTAIzJC4efK+BxccSBcz7aKKSFoiFMIGV2pIIgmv1snzHw7P6pPPgfpcp8519PgHCRWFGP9IUbeCVCukLoE8k0u3IqSPyEnNUiUVgTb1iy9OBdoyU4MagA+Of1jJSgpLExImsb7M/GdBO0h1C9WtyppVFzhYgWMBM0SwwQxF/unGoEwAfJUqDv/M6k89pxJmkyTMEEgTKf6J0qBlvUqFzFANUqWrcLdCxKAIvGr1n3LPbAskPKf6hdMH/0FHIHSuAeldgzg1U1UJ3YrmlFNsdU9Ngb5x8geDZE0I1/f+dY9XiBMyNaFvGmjgGxvAsEWgPwSywQkzulmBqm66YacXUv7J55+SN4nWoE2ESWJmac961U56BOpWoCQoG4iRcPA0kbJ076oXJF3+4WGgp/9huF9w2HX/khUeUmFF1ab/6RrhvgDWqhlnqUpl6YHQBsnhgXABiRWt201IirJJnXKsu0kVgKry/oHBYMDPmiIrVAIXyJ5/Lt5KmYEecFyrwumTwaC9UwWpg4EwN9xikJQA6YHNQxd99JAiSch0g67JUqBHBPKGdCS/8PufCwT6u69QMs37HzwSWt0sIEAfiAX0fh9oCYHKAAmA3sWe6gPYQyLeIDUEAnsqzZ90PnqtBuDeq2NCqnyqRwD5/i77EsL0fK8ERFIL9mGfwKC+47cfvosbySp90ce////N5SAH/1BBD3ZRi1qA4A1vAMAbAqAeOEzJVARQQEJMAJ8KjgUOCTrL/ACI/yT7RMNNH7TVMkKCKv65Z2+7yxQQivAPCZCwK08QSPYCFwuDAEAgOqxGSMoxEExQpRzlmMII3HAILminPDpMSAyfxMHbdcV7o2PAP6pIKueNUIaiS6FbAmArxXWFhSGJIgAP8Z4MDqQHjJuEF/7xw4GELyHlmMRA6iiQO/4jj1PZI+PK4YUpsOACJRgB8mj3D6ycqQRbZGRCuthISEYSf4BLYw/geB866hEkl9wkVdwYSEok4h+HKMATCuAk5Unyfgp4xT8KlqkNtNIs+vsHB1V5S0m6wVZe4OR9JgGAHZhyIGwwiAv6kkpcfi93A2mdk0zxD2L+owvo0c7/TBVGbv+8KJnb9EodAdDDf7jxSSb8hx9DAs4oJHEDxuRmO915vgeF8T31GMg1GuGod9ZwIIk8kzi14sZlgPM9wvsHQT15yR4MIJrHzGdDDcbO85nPVqgTCEVJmLeLyU4gpxznQMoxghn8Y3AGNcgfqzGJHjJxIIwTSC8H4kYvKOMY1TjGD//4x3AOZBksFUhNa5oQC/iBDYvQTlMcelSkJtWaCVlkC7wSixG88Y08Tcgy4Fi9f+RipDnNij/HsowgclUZJrSqFzAxibMCgIl7++JA9CfRBsEhDUoYQDXlRrpxPImeSg1c5P6xTL5qRZ6QNKRW1tIDFgzOo1OB4xSM8Q9LjMD/pUjyakkfUI7Lgi6zJRXIA1h62Z0ORAACIAACjBpY+mgAtZBbLals+L810KIHlqQKSUUK2U5I9pKTpQo5W+qWyVJVqgUd3FaF+49YEOBcrWWurRQA2IT9wwLw2+aUatVcg8w1qow7LlVmkIv58JYr1ajGEOfoFWU8YAqK3W1n2WuQ46p0udhtJPTOl0b6RO2DAPCf/S44lcEKTnAzmAFvFauVcgh0CrGYwRRs60MiBsMQhhiBgxcr0hFI9rwG4eU/elgNqXAFmfQ1mOLsKxA/cIHEjTTVGtRGugCTqoheaax612sQHBoiGDsQyBSI2FIilmCkUwipQNBgCUP4OKpR/y3ihIOABiYzFiQ0iGDiQtK1FZfYygkRJVcqMRCn2u8N8KmcSgWC0SwnpHVhlAALliCDL/thilQ58D+AkBDGabage9ZzSA48xKi2Yr1RFUgwgPFbzfqYyIZ4wy7eEAyDoIEKBhhCFUbAh3+g4R8jMMQ/qPCPFGTlwTv4UVTGjIJHjuWK8EFcV4ipHQ7Yz68JmdIYuVnY+/Q3zQKZJlckcAFKPIEPoWwBL7jgBz/wwg/GqEIs+NCKJ8ygBFjVijJUwAIV/JCniZ6CIXC4g1h0OtOeRoMk/lGsfxhDDdw2xoTRoGmBVMHTwBiCuf8BhiEkRNL/kEQfbtGEIVBYsTOunv/wWBrIcugwEPPRERxiHLpWZ+WKrwbgHEJS60n5YHPIm96uuaeDN/+jBIloAbb/MUAVJITaLGhFyg1S5x5vepErdfAIYlGFfxtjBBI2siTq/Q+HDOSxNkbDhCNNBZ83QSB96IMtyHCUgUi63rcQyC36IAlJBGPQQTBAEGYwAkcIhNDVK/JAwGGqVvfO42sfC/EIjSQzd+WMPZhoJNr6jzt8kAu8IB5WqT0QwTD8HzOIBcw724NcCAQYt5BEIaD+B3MPYepUB0kI+mDpJhukCpSWxC0oP5AFOKMPSgcGMAxQiJD1QSC26EMIxnALcWT60ymQNJQHnfhLf1og5IAD/x7/PpZqQojtzB1BEAOATwBlydZaScBAeg0g04V1cnofCB+moAasksFpvqhCIAbXCUpA+sDVWy/OQ2AQOkTnNrgBSTjM0IRf+GIMO5CwJIRGdab3YQEx0K9A8tCLgVCJf2CH9rMD2Ds0ZMgCYKgCKqCwj+o0NAgCHYuqWAgEdMCy5Ru+1pIlDQSereCfMsqUWbCifzi2feCFXMgwTku8bfgHMFG6fxA3oxO8HmOBZ0CHGNgRr8AFVbEDO2CFWlmABXiaH+RBt7Ecr9iEf9gEcPgFrGsCMLiCFDCAf5DAYJgBS/A0A8gAKjSEBqQCKhCHMagV+7iHu+vA1fqvhODAgYiA//rRQI3iiiM0GC6YhTr8BxQcghTgghTIgBTYhwzww6CrOn4TiCBIiMFRgylQAWMgBzIBiUf4Bh+kijnkiv6jCiz7hxjIDxuAPMnzNN0LAirIAHnww64zhEDYAUZEhzVoAHpqgNcxi0VIiIUymFhDw/t4Plx0K0biAl/8Bz4gNE4LgkPLinzztAz4hwxIvB7bOao7lq3AhUpMiKapFV3YHrewAx74GMYbgq7ruiAIAnlIAXMzgFC0vgcIBGM4AY0RCCK5M4GgrqkQjIF4JrdQrb64xV08i1JICAdwi1rgHgtgOw/6h1vkgn2ghBGonhGwhEMUCN1LCIwAg6OgNCoYg/8Q+Ld/6L5AeAZ3MIhMHIjrAolpNAhW4EEkvIso7Lp/oEJ5MAAqrEKQ0Lr1MgYUaEV7Gch93EmHkpG7eKGsaKbR4QA/mIHqMQQDKEavODRJGEJNHINRGIOq4QEewMb3CEmq4AFtNAhJMIAU0MOXNMSp0D0qaLDBCQRySIMGuBeV40lJAspJuYT3WKS3y6cwGjGBSDUH0MV85AIG8IMU/C4DyMKYTIhDi8isOEJVscrAwYWmqRpDLMyxOETbewBGpIFs6AEBckvOfJK7sYvp+x5lgEcA4oARrAIKiIVYsATJ7IqHdJLrYkzSeTLsUwM3MAY3E4gBsoItUrHOHItSEIX/30wI0rSfKyIEJciFWOiEFECyzWtNkFDKqRjEoxJFmhwBSmiFEliCEhggvtgW7mFGgaAhRgKbM+xAjuKofbzFD6AFciCAYDCA8EMDmIxJ6ByI12xNxFQqNBg0SmCCMqhLd/oySXIf0hmVfZTLF1pQ0SFPrqCBN4g9SghGLJTMUAOJpCw9cQCG2PsHcTA3SWCOSXGCf5BOw3lI2/uHJxikfwir4USS8ySVvBpOHQKC8nhDwBFKregP2PiHZ2g2QmsFS7jQqaBCccCAU3iHdzCUnjEYQxEIeqAHCiCDIXhNEyWVr/uoVgiEAGDLF72PGOWLBnmxuwhNJHFQg6ClLw0J/3VMBBYoMuaEznybwhQQBwpoBtIYnZ5xBTK40sChgicbgR0ooiiIA4xb0y+tnfQQLUQ1iAHIi/nIBUogpH9gAdbMihQABgrwGdF5UlfAAT99DyIlUqoIx0+bgUCohkAYgSgIhFITCCwgIUX1it+binYwHCvwTsDRyYHYg0OCj1TwUqDKRfpggoTQJSe51TOxgECQVEILhiH9h2MENdxgBBIQAYE4v8DZhKRRQvt5TSqwvUkoBxUgua2QBY2DnVm1lQPoQFN4JnvcCl9dVxJTrXR9EroTiEPIhSIDhuiwAR1kH5v5B39A0A8quk2zqRHIBQKggTWAg3GxH19t1G2CBv9bea3xEggviLvAUYGBFIeO8IoYiJ54QZL71IppTQgqhDcje7evWy8iYoFcYIBhGIZ/0Lh7xcf/qRGBGDP40EmW8oN2KoCO8zihVSV5M4sfiIGk6cyIDFeoDcdgCAYVXNhVmId/0FnftJ+B5LH74FWBCLNtKgC6A1sA+q9/fA96NQuV8oKNpVj6SIFRHQhSpYpkNIiUDYlPE8VwhMnm7AQCI7BW4ARRkIUW6DK49YrivA+Xm4pZ/Id4HQtjRRI1hB1wqqwPGln60FxNHIiR5VzSuVu+mNa6NQhRrEK/9Uqv5AXAvcJc4IUWiIUeSbXE+YFk+QefnArEURieXNwzidf/yN2KUyJQn2Uf8TwLfbmlCABdJGFerYgahhGTTJnTkChduu0KKqxP1dVDP0yBViCwWMiFQ8gGNBOIaWiACJCDWtSKe5BNUtHZxAWQC6rc0WkEXfugpp0UW0A3MDAIRhCIT/gHlgFg0RHdrsiAfMvbqTA9r+xDB0bgFOADZyuBXHgGNWlFjdGYZrgBYtoAg2AA0yKAQPAFRxMdZRWIe70foGzcs9BVRqLf89kjgZAos9gBHltb+sgWxAAcIwCJT+jhlgkdAz6TmJRbPwxEJObCYGCwVsiFMRAABtqFRkgDONCEIeAEBuCCROBXFgApPiCEbEiDYiherUjh/yleJoLL/9ERJ3gs2heVYfSYgVbIp3eoB2dQhAC+t49R0kfYBCfIYyP4hE/oBmwoSUmSW+5F4izIgCxIASrAtFZISD6YZGAMqRngg0vO5O9NBDfwWoNZ30zZC5+VHTe+jypatRUTWkwQqEwBHcw1C0wbnQhYgFmmD2wAiUDOkUd4B4K1hx/4AwK0hW3h5UzJAic5xq904EXOgiwoRXngBTR4Nl74h6nlA0PoBEuwBEAERO+lghPMisQ7XvSAKFsx24GYuS+Fh7EQKE/exabN37vAhkfwh4FwBnt2hhhQmHfwh2aiZ1IxZpCACPgA6IHItyMeAmMmaGPOgAbkg1zYB2bIgG3Igv+JZuZtGIJtCD6D0WiDMectgoq9iJ8uKIUu4EuvcFHK0iTmO5MQgyR/fodCRhJjlgeBGOKBEOh/wOmtwIh/IGiDSIEepls/XGZjFugjOAJ5sIRO6ARD4AV+kIdCEIOhwOJ/mEVUthVTcIHg9ThvsCj3EOfRYSJwwqHvCVOz8IMX+IIveAM8gIodWIILMCVFbVeBkF6DAE/uuWX0SIaEoOmByAIxCImP4OmuCOytYORkZOYsOOqjbgPG5gcUNIRckGxe0AZOYIZb5AQEqIQdWCAL2IHPHlSBINCtIGOQqCKO3gqP5iuvNpzURg+OPRMgWAbQaW0n8UU5UAG2/gIA2AX/AcCEHHiCFb0ALjCBeJgHKDgUQMkyjOCHu+ANjzAInd6Ko6YIizgCZLAIMWAGXgiCJu6EXAA/SpjmE6QE1RyBHsgwxLOEFmjvFrA4rgiiOEzcx0UANBygy5qKwjEmcr6PXWhrAQAAFYiFEniCVpgAE3gFBU9u6RWTutk1wqYPh5jwjPAIZNCNNriINuCHDd/wbciAE+QFKrAESvgHbMZmSxCHPww/StgHfdSKBVrTFyvIvpiPvcDRd5JHgehv9LBvEpwKYwDMXCA5XuAFSijxVmiFTmgFcYgOuwYJeI6eKH8nw/6ICheIjxhsDb9wMcju7BaDbeAHiU6BXIhlrUBp/6rYWq2Arq81CDO/D3q8i+sBEBAI6dUyptwJBQ/wikWaPgtAVoFAgPnxnigAgbVeawDogSKf42drBUpgaj4IBj6gTubWivU7EyuHAGQggY3wiYHoDd7gjQtHhuyGjm2Ign9oZ4P4xxn9BzakCvv2cYNp6al48/tYivh9D/4OifUxiNki8Fjw2DsYgAFAgAHggmMfAD+IghcAgf/2bQCwgC6egfF+tmBIciXvQwEEELzmppANHWQ4AuhYCVDIg1XAgUBYoBgfszfIu6lIW4F4LPuh9X+gQVuRg4Roq72531vC2KwoZfcA+ITYc7NgARawABDoATkYgFCABmhgA07wxf/bvANjYDZLGAIUfDZrV/J9kIeJnu6A/Z5uN5hv54vbuHSQyPKEsHKq+HDmoLc/5IJtYI5cyAVjwCE0DQmCz/X7APS+QFb4th+y/od8dQ/SBAE8CARxkAM/sO8iL3KJ5oXBBIZsHm9eAESBMGaH8GmuGPkzyY9sEYgdNggxCXkA4YhPBxCWTwiUNwiSgAASgHvfmPtVYAZxeN0hCOfhOy0AQgFUby0cEnj6qAKjkgMiQIBQ2AanZj+exogjAGiC9mut/we/Vu7QEZok1JGu4IkMx3KDaPt/6IjboAMoAAWf8PSeOJP16wihiHuhkHsIGMchEAcFovepSNreyX3Tdij/vnfU7/EEgSj60bGLRvCF+b6PvHsGABmzyjleOWiKhdM+6HBugTDsnD6CbXACMriBJliBJNAETcgEkwkBJxiP+AmH1RABRmAECPjfqWh792e/94/7rNgIKJiO0P+Hbb+P1gcIEgIHkkB2BUGVN292ocDz78u/iBIn/gtFMaLDixo3cuzo8SPIkBRviAQkUqSvfyBOnhQhEsW/SBFNsuQoIOUuATV3eiQQkQaNf7sCpCREgMu2VR5wCLvorNk/qDyn/qvB0pWIQv+y/Dsi5giyf/z+tYl4BAIoOqv+hT1JkAQogf/yzI2YFoKkKkO2/aNDJyKJPCQi0qUrcTAEEhBW/yVurFhgnjx0Qm0TJ0dizn86/6WkqtGn59CiR58McOlfxoiNYooMRHrjh4tBX9OufdJZRNznItL7Nygi1n4sYYkk/q93jRURjWuERa3flSMTj4AFK6YNsjZlyYLKIw5H942DOcYtDzfwecGg0v7Nw+hKKA8i4Hu4UjmXOAIEsFSJEmjXUBNFUQVooIX0zGix2bbgR1gwGFE0HcVxUS0SBaWERC9Y+CCHHXpWYUSX7HKRgtS40lRUFfT2G4v9uPJbTcTBAssKNdCjhx7NQHXODx0lkdxGGJxByBVrmdXGddlp1wYETC6GDChXPHPTJShEIQ5fadX1zyqM/OMlRenBxf+eWleIQ0ZECJzkzT9sxlTMPxjupKGHddopUhqvuXnRGf8EdUJEiPwkURgMWvPPNYDQcudOMol2SZ9yTnQDDppIJFUFwrhSVaYTKUfRICvUWMM6FUQkFW4R7VbTORX8OAg11GAgKRb8UeDEKoIVhAwyEPjaq69MXpFHAv88Q8MlvuyiBApnoMCssyjsQoMSWBBCwbWEYIAFOSnVcto/l2DwUkQBMHrugoH0WdsWhWoUYZ06gLRFHeeymQ1NH3XGYaKHTvQLSIvuO6lEJNUghTArhKNHBaZ2tFuq/5yzqsS57XZOxFRVoFzCylVJjkRbSGTDyP+QcQMZGIzhy8r/mAv/J0UYyivviB11W9O66IIkREQO6hySpD/TVguIgAr9kb8nVVhMheBKJK/QtMDckRmu1OBwxVRRfOo/GXMkVVQareBKqUn8w/M/9dY7EQUcAVpLMVL/syiI/8D0kw5AibTo0R/2vVEqf2vUwD+EUwTHRfB6pkqH8hbDOEU0TaizFCchPhEkgoI02z9bVG0Viv9gTdU6H0UcMcQdiSpMpytgcALnVMGZzUdG2xb7SSfwPdqitPdNC+MAqxJ4oFRVHtoaFBn+UfIgaR4R5HdGIPhEmfxjKUh2aMQNNx6pogotiCzwolUarRN6baVfNLpHwtQQzvmlu+qKyGj/g0RoqgAs/9H+1MvGUvk2sjvRCA8dFIGc7+xHEQNKhHjEEw0kTgCJOi1PJA8cDf4iokA7RY9DcGheNNYwDZDoQhepiMMvyMAIkplNIt2ISFPQxxMZRgRr+IuhRkylPor8KAk7LN0KqLECGnrmef77CDgmR5HKYe8fghBZTaD2j+lJpDccEVTg0JGvuU3xBAv4hxT/cYITQO6CtWGFRKh4xIigMSK66AjYRkO87lEkT2uMSPKa9w84XE4ja7ADHLQXEUX8QxGEvKNnkuCKGlXFdhKx3wY5YkaeKBEk+9MfIkdDx1SgY3iIUONGpNFGjQiKih08yShBeUdcSEMjp8AcD04ihVdOcf8iE5oQHVlRQqoo8Y3/GCVtKniR5n1RIoe0gRPCsZEWSoQRiujGOsxWuk3YSRjW/Ag1FZEMdqwgCWajwCkmWEyJjJOEk9xILDVyzo7QcifAFA3xevSP452knReJwxwpMkGJQMKX/4gGLiaii3ROJHAPpGdEyimREe5EjxO5B2mEGaFHhGSUfQzJKfzxj1cyEEKeaeU/TigRxXnmoiBZABgUEYKI/IGlyfzHCz3ihGTkoxeMIEU+/pGMf7DjItSc5muSY4YaMHMiZthpTv/Ri3H040f/sJ7ooCLPk0zunQ3cqEYlEssJmbCSZ2RFOkEqETvWZJL7nCpPiOdVbqSCB6r/lEj3WhmNR/SxjWh8ZSre6M9M8lUCfBWcRRQQGi2EhKzCvAgn/gEAlsyBNCX4xxKKMJEAkJV6XIjICxz6181ydioCEMCeLtKDzpIWJIT9R2WnIlmdLeEfj62jaLogmglEZAK0BUkOSqtbW/rPXP8wyWoiQkeN3I2vifWIV/+hAtKgojab0UhqO6ImjkjArxMxBUWKtRPrlgGyQFhsakLjAOPV9rYnae1pdyuRSmz2sHdaLEWeGxLfqre+FwktS+T7D0f84wFT+EhzOaLZiDC0iPZFV0AXNI4DCw0iDJYI31jwDxk8uMIWvvCCaGteDIOEThNx72bT21mTaoTEGskt/4cGrFva+qG4DFIxh0VCuOB6iMYeotMdYjyaANc4Dg5t21RgUJvRikSPLTjaAM7lqIkUQMccATGDbMwhIDhZcHBAx90eO4Me9IBOUViua0CAAl/4Ah3oqMUN1tLYxuLWIxZhkEn9QJENV7nOEmHA0XwL30zu2c4SCTCbO3KIfww6EFGQyA6qERFFR2Sxk/jHoxfb53+8wQJR6METDsEFbShgLR7QSGv/YV3akDQiK3nyROiMrsvcKWlVnu7fIpHcKdf5CaPBM0WanIsnjADSF3H0P7wgEWGz5NERWa6t37ADdEkYsiX2H64ZtQYY+7naE1ltTYQs5DV2IDSoECxF2P97bGUYOyLH+AejPaLoc6e7I+X2dUQeu4R5/wPFHHqttYs8Ed/lrh4TMXG+Bbe86P7DwzWhcPE4/GY1sfe/kD73nZbxj3IM+9FLeEIZQh0SF1Clu90NeJ2aB4dxgZy0kxYJwvmaCNGEghexUMZFhC1xYv9D4h9pd7CHLZF0C5vmFJnEJLwwAhaUwNYRsbWCJILdmgzM2SV/OtSjTprlwvs16VY0zYVdjaBLhOIb8fo/lKGCXFBi0BJZxHGpgm+pvybAJClt2tku94lQ5uVTWbe6J47uiU9C0eXoO9/B3pG/b/0fanhCkyPChtF8fO0iSfLcJwJuDnH8HyaoiZQjUvn/yHMe24L/iLE/e3KdR8TnGjF9zHWu6MIrIxa5+Edi474Tx3O+zkuOyCKuy1er1v6O9P38a8AO/IlMwQ/a2HzvL0L1amvgI7fHffKjHxLTQ1xo7e7BZRf/j9xLXzNbpHZ9DxCRBXvk+aPRI5TXSJNIeMP8DF45h/6+EazvvNyAZ4nPZZ7zmce8HMR+9A4kwuK5wNKJhKBoHEtEG2ctX501X/clDiCsRnC5X32xV7fBn230nP/5388Fm9dBHCb03btthMRtoM/xHwpqxAP8n0R8wGVxH098XE1A3gP+FfIJjfmlX21QoM6EQqDthLhJBBF0hIPVxAP8wwiMQDkMn/9V/wMA9JkAAADXfYTNccQDLMMRXuFECN/eacY/uME2wCCHXFYNlqEZRsTksUS3dRtIREGzdUQVruAUzMA/sID/VeGwHYMX/J3WRcQIdgTNRZpi+ZoIhmDhodsksJsfSgR8EQKscYiqfcR4nSElRh9hIaBH6MRyeR3Mwdzw9RcS8kEuxMISHqG6/SFITILgQRwA6MRnfVYABEAkyCItNoItFkMkFIONFQMhcMJ08Z7OlAIiOYFETGIlHmOH0NESjFom/kMgxMIUmGJEUBzMUQSxzUAsWIISgh3qhQbFfaPeTeMe9lzNNVpEbAZ8xWIkREIjAEIapEEtEAACiKGOBQ0ydv8WfZ2hMoYEIAjADsTCDiiDNHZd6kUEFRgCxQ1kzpEGOIpjRDzAA8CcKUJkRNgcB+IhJixWAAhAAKAAESQWQUkfNYlC7fGY1M3agw3hPzDUatwBkX3EQB7kFPjcJ1KFFwxkFdLcES5DOZii1xFbFkoEHkZEFODAP4Tkg0XiPW6ESS6lermhw3HE541AJ2hjTy7kVNxkSPhkf0mcQlJEQmoEK/4DJhwCBeyTU0YftnUfG27WLwBkTVajRChDOcTCPwRDVFZkTchlTdTkRMilNH6lREQBIaTl06HCHDTlRlAZlYXEtv3N2kTENYAE+E2ESpYWCyybSCzhPxjCCGgmS1D/ZDnwJEh8XlhCJBOGI0Fu4UW4BspFRMoZ5oElgDlwxFoeWPLUzRmWw7JBo2gomkIKpjX2ZDn81wN83hEKZETkpWr63C40XUfEpmweGGK+hjH8Q+JZ2T8kz9REHcw1Jkgc4QzsQESqpkh4QSum2wiogUgc5z8GQzhSGcxFI3GGnX2OxqH9Q3cxgWtN50dkJ/WA25sFHEciknYNzrk8wAgw4NdRhCf2lzR63QhQJGtOxBEuYa/9AyUYAlhO3BTwwQxE43+Z5kagQ2X650csTxihKG1sUe315HoOHkHK5ecFAh3yQTRaaNgdpzI4nH/R4T+gARUEQ3FGZXHOgCEYAnwu/+dFSKMXnNsb+ALAsShLONKF6Zd68WBENEAcaOm5gBgC+stkbgR/gUQ0qgB7TmSHTuNDTkESmuIcRkQuKCEoPuRxPsAM9Jp/jQAaRAQaCGkn7ICbGt4/7MAIGAIV/EOisilHeIGwvcE/7BWVnoR7YaB98aW15SOHvIJEyNZFVFBKSMASdNeR/UOSDYAcyBnsFKpEiBhFmCIQ+KR/aYRx2uc37sAMBIMSDupdokEVqAB5Uhx9lsMI8MEICMAbTEErLOmfAsMQWIKh8oEhBMIcdgIaGEAGAAMSasSDTsSygUOkhhQ6+EIgCIEO2sm58hWPKSaj+MA/tMO7TqrOeCqqUf+EBJTA2snZRKyoGrBnmc4lt/6lfXar3kHkHHqmm/5pkGprFUwBNbbpCATDeO5CMHCoRFSBJORFE/SawsKnkOYFmXJlNU6CZtZMRARCIPhCunoI4azsPyweB/hPGm7EiUpfzVYZvYJESlRCC/AsL3BBC3CBH7SAHyRZIDyDMUyBCuQAH7AAe6pgRFDZFIgdEHQiwNKn0nqonwapRCRqouKlRBznFFQshwYDGlisojrrP/RBEwzBRaCB2kYEMCxpFqrBEjztReTADsCXa4aU4ZisztxsGcIrvIpflqZlZ1BCK4xAbuXADPABH8TCE/DBE7BALMzADFgBe47Av3LEFAD/wQzYm0TQ5w4YAyEYg6BKa2cGQxX4qiRERCGQQS4YJ4ZK69lShJAWAjJoRSGAwRBUQRVcrF40wS38wy1IAhX0miM4rChmKEWoQQ543X+9wRiogsuuEXbRY98kptQJgKvJK0gIWQkwgcsxKKE63H+pAQvwwT9MQXp1btgmoWoeJ7EGwy3cQjDg6j8Eb5BSweu2RR8EA+r216AmKddGRBU4axNEBNuSwRC4rUHCrSQscPGGwB8AwwgEwo925gj8F3+Z4gjk6V064z8swPVmkgKC70kUoQrvRCKgKd6mb/tGRL/+gxXQcEco6AyogaxOgTFUgTvcr64awp9WgQFMsESQ/0EICPEO8CaScqjXKuo//G7xwlQfXHETGEDwfuwQ3C8D30IWh+jY8oIBoAHYOoIaYG60toJEBMMuCO4acYAcH1ECFAsqHGgL942NjZ7gHFkL8MJ6Qi/xne8/5MLydfAM/yuVscDrGUMSuuYt9MH93oIED8ECU0QIXDH+CuoMdELXwu0/SEIVM/AVS7IklDEVKHDxVnEf/EMTSEIwmK0BpEAQmPEUROOhti8dLukzLEDznPBHGEger5HeRoSX2gkm7mAjOAqWIpIfzIAK/Bdz8gI5oMB1RkQsGGvUSoTUvh7+SgIpSEQyJAMjMMLuhvJErNTaanIHwyeHAu8Rvy4Dw//UF9lBDIxBxoayJbuyRNhCCIxBDOzC66byECTq2d7ywXpmK3SCIQAvOvQRMFOE9g5zJi1bM/MEsQlAJExp3xzzGnHBnE7EacUAOChB3/5DK0RlVCqoMYyyR8TDRYBBIIwByh4qKE8wK/fBGAD0PygTFEDBP+TDX/zFROxURMSAHeCzERcCBJ9thgYDQ/fpP7hcIGQDRHvGRFP0HUFqh8DxucildEpERNOGvvLC5E6EOEQqwFyzxTrvPxDW8o5A8KqzSOAGEoDDLxxt8JLDTv+DO/SBO4xCDPCAIIlzQUTEFUyE1/xBDCCIs/LKolJBIBiqQfJCEOxAIDwyCSO1RHT/p1Zv1uV99oOQ4T9EWy7wQUqj7DVPBIJsLSK773L6sGu4A5oYr0YktkTUwxrgAi7wwC/8gi7AASuMQmAvQAz8gx28kShNBExzBEPZQAjY8/BqxRC8riF0gvMacQoYgEQoqQBXwRh8Q2eLNmfl7BlCHDMqz0Qkc228Hq5NAAP8LC9QghokoSdbgkTcc0QEA/tyqCe7xhSoAX8BwQgYgy9Iakc4jF4h93K/ES4Id4QoTmGLBBKsQQy4w0qxwx8MATBQgYfzqYdTQQpst5CigSXwQgqEd33Nwp2RN/RIH3yBZ0dwdG1cFotzAS/kQiBULH4bQBBw9z/g9hI3Af9yhBa4/6kxgIMuFHZya4Q8KfdIJdhGTHhNOMMoDFLbIq+HC6miGoAYZMA/ZEAGWMJ4GgMKrEEDjLXQsPg/xKy8voJ5T4RX+xn7uUxIONQbvkZ+RkQBlCoXcMEscAEzMEMG5IIldAKiG4AlcHdb/EMILHCHGySita/D9sAz9PVf/UHbaisV1HKXg7lE1PKEqkEP+MK0dTYmdEg7kN8/OCBPcABtkTaLxjn/9J6mUoSVHg2gA7rLPW3E4reiLqpEvDIE/0MQpAAES/MUBAJ4b4SUOzuH+JMtbHoQGCQVGIA8RLpEdIIYjwA56AKUuWpHZG9IuKuL8wStCwq+ggRF/cP3cshj9v/NKQnOn+eCGtxwZ+K3tmrE8f4Dd++7tuJ3kY7AM4CMVlEFgoeGpm94RARBECRqBgB513ZCSv+XMdAAmkdENqS6RODtRsiem5+7bUyiMWoE7Y0IROc6g8iAG/xDLJzaTtBgaKR339xWoFMCinWytu67sUsEBIRFFqfAPyiw8UrC67WvXF9Ewk/5RpQQK+CCLtWE9oABPxd02op5w0vxomL3mXrCL6T5P/gO/D7IMIj8RwhjRJR8SOCX2XsEjodaMARBh3O3xE8Ed0PAP0BAFvzuP4yB8B4tOQB3LCElRVB5R+jR0l8ED4BrmBQC8gJDCmSBtmsEFYToEY7AGcAB4Rj/kMe3/VKG9VT4QWHqmJrgeIYaArB3BDBUu7FTwRA4/mDHAHF3g3H/whjwAC44+LNHRGEn/r8lmO93hCIs8HangDwYgIf3vEYEgWcumw+feQMwTud7PvVziBLgW3eF10XQek1wgI1zwXpS5Y+zPs9PRLVzN+tP8USAQwz8AmGjkS4Bo4f4U/ECAy+EuTyIQ/J/BEMDxJQpjqZE+dUAnYUc/7T8Y+gQYkSJEylWtHgRY0aNGzl29PgRZMh/b/5FE3kSZUqQL1R+5OBwwoBYI0ZQsnQR2EUyEO3g+sfKDiuHQVMS9WiHh8QgwFIAo0Ilo4F/QaCOmOJQRZQ46CI2bPkV/2xYsWPJVgTxD05ZtWKBUGxgscRaBhEn+Jk5IshNvR2DOHzmUOg/o7oCr6VoR5dSiH0xQg0i9R+aGVenxELxS4XDhYY5d/YM8apnByBNqoxr0dpnjpj+KcNY76SJlgQ+xJrKa+piiFQMMBZphyNSslBF9qUyQo2jHLHO5FiSY7Pqj2wgKtm4R3p2sKO1ayzW/aJriMvAY5xAActMSzcj5vT9D3J58AagorGqZsQHFqetRJdfkY2XQpKgrHH+OxDBBOUzBSIMPMllBCpwQ+Mf9yIyICeHciJOQcOIM0QNNbR4IpcSTjsJuH8ySxA7w9rp8KRSYKxIBohqzI61GSkihP+GKv4xZD0+qNArJ2DYo+i9InVUibgg7JtCjVYoWaKEJZYQ0aE4luwoF85e3BJMkAoIE0EuPqAFg8h4sWSETtiDCsOO6JOETJQ6sWqKCyopYwmJtOyolhmfqFPBUwg9NLuXCGiEnFyAvBMNSwwQB6IMK6z0H6gcc4g++uZziEOxoLrzqhIo+efEABBdVccu5GPp0CKyWwMFjQSsJZBccrEERD4ktVQqSx16DL6+LFRS2K984mGUiEL9LAirUMWuT1athSgNtMrjzqG3rh3LEYmAaAsiWWdE4B8UQDAml1hm+GeGTgzAjVKKgq1CHAooqIKCJvrVNxwKbqAzLHauwBT/ovg6C6KTYASyYsoVv51YVVYjEOkJPmyb8Q0BBJhIVnN1BMQhEO6ogiYr/mklBdw4lQgycapYIJpHTtFDj4tCEGmLibaooYYVVnCFDDKONOwmxoKYYYRyouSjGlXTmpjqqjsi0GrOTqyIC4l2OWSmJWbwFbdkJ3Lnh2nIAiMiJzDS5IaFJ+rLEIEeKIEFAeJYI2syG+l7rr5V02AsPNygZIQ+Z7DEZfgwzVAcDH545z9YcABGYbmnaniKclQwphg4vBU8zIpVCsD0JS9wiImJaCEdI8LJsiCKXPgQu01LmnJo9396lwQDKZrJuTyiwTMusqZ3COSfvUeHXaUwrNsS/wCQRpjoxowYDImFS6CXD4Rcc1kicV9jrkicJoT5bwUyJFFSuyAYmyGQat4IJJBs0qzohO/Bqzg0B1odWQY1QId4zyG7+McX/AeSbIUkFodgwQysEK8UZC5h/wAePSKiic+sI2f0cIU4zKadUd1pB9X4B/4Q2ECN+OAfX/qH7GQXlh2o7B/+cSFE8LDDz1ggELzgw/XgZQAMahBDQ7DBgZxQL+lgMGkOQeEk/kFERLWITKnr0AANmJFFcEJAFKnYE7row+68AAQfyMUMFBcEl6XAIRCYiDO0U4F/pAIiWyDYWODIu42850leUNEheNECi+CgQyzgTA3NiBFTLCIkrf+r06A4QsXYdaYHtrveCPgAjCvkgRHhoAgPYlAeHuAxTIagXzUmsYNYJIILscDjGr7TSFtyJHD/2F5GWuGQMm4Ja2TRgAzHYoF/xIJN/6CUKJckjHWg0jBH/GNEmLaDf3hBGSMwBgrQ8R2JVWQYZAoiRoj5FS3eknVfkc2hGKkW2uGrEBG5GEV+IB+TbAJMdApVMIKBnHLsYAcjiMUTbBPOiMBQIp6A5oEe+MCPtFMi1uTIOVnFiQYm4h8dAIkl9yYdFVgAVhRYgEfmic6QoAENwUBDKyYjEDUsgRLbiMc8/kFTmh4gTB8TC2tyZFKfYoRkHo1IKf9BR4wQtSKP+On/RlCK0jsFYgo0MdUqaApRGEnUIy8qp0WisFTtJOAVq9mIa/zAKuYh8h808EgMkPoRSPi0qSh9ipOYVtdWcOIVPhAFTrck0S5xZKsUEY/VjAmmdXILLLDyiCBhVFKf9vEjQ4CIZC+iKSpQpTe9kYxdmZEOH7iqElYLbEWwOjFKhmmdHWKsD98qEXAoCI6QBQllOTLXxxggBbwaAQVnkItVrMKrZtxld9aZ2v+sdkZSUMtrEyTbiDg3LJqSnxEvmNtOzAC7MzhVaNWCxeDiUiVlZYMpwEgdjpw2LPBIgHz+VqdSxsCxYkkFD14LjqQYhrYdge5Xpotb3KYgBUEIBnZH/5AL3PjCIfegyDTWAAe+veYfCoaId7+LEXSFhQ0bAAl3VbJeiHi4wkf9B3zhS5b5QuS+qLxvA29L3f+m4Lq7jQUvAuHQiTQgAhT4hxw4kpi/hphcFMnlhcUSRo4wIYAtASt4ABEJRMVgpGNBpT8cAg4qQ4S5KJYINirQLIhQDiNL9Mx+k9UXI1I3BRlIwRDWlF0+5EKto3tLAxpQj1Tw2KL/gCREoPm8TErHQCGWyJ61YwJDyyeolgRT/1TTjYwogm0UUcRJMvCP/E5EspXGiKYv8p5/SOrMAAawmlNABWOMjQ9V+EVa+EZnV//gBnveACfYUGsikIMcv8hWUC3iWf/DGFQkbdGpoKmWaOQuiY50jC9YSPGJfzS7Ikb4D6cxPVlLW/tlDtHnhUK95jRnIAO8oMLYZtCKXByEzqJzNSRuwCBOaOMf2mDGNngRC2NEwRcksZpOh/2fBxD7I7w+9oz6t+yyfMLZEfkEKaZ97Y/sN1i6kcqLvw3uDDQMu3x4hi7QcQk81EIXdI7ADV7CAW1wQYgZNwaCFXgWi5QChl8KdIdUGBGd6jAkQf6IIL0CcNVINIAUtpYijOBsaTM84YyQSC8+YYRJPzvhYJImxS0Obl50Al7/4MUHotADY2gzFlUgAC8oQYlYuGsGEyww6LKl77KYtzMk6eFXdG5LeED/JKxWa8vWJvaNf2BjDJF2SB++8Q3AO0Ha/zBC0buRFGz8A5+sQvOoqz4EAxgiGP+gBC/axYfsfh67ZZiB6LGbCxW8wZpuxwhCdcRAa/awh0UIpnx67vO19FRWBFLkxJT6j0fgIhxs+8M/bHFfe3zD0dIm+uLHEANcvOPKX7l0S/qYgj1KQtQVz0AWwG2JXmqeF+V+F7k/z4dOrDEYuWBBOTyTZ8PIyuXVa0kRYFV3PRN5AmLNGhEiAlDb/yMComxtiM/pxuAbKOfxviEEPuHpFMHRes9aqO7buI/7liYYWmEfKGHABszzLpBx9uHqZoAXMMohVE8+KKW06mQR8m+s/0iHBA3j36jmFxxiAWYQLO5hHRzCFowADHbGIZQKGx7BGRytLLKgIoyQLP5rCNIsBbJgCCgwC2DMEPiAEkBQ63ih6iyOFwyBF5jhx/5PJHgMDJeqpAwOJCiHcpzBFhThDxQhBIzqH9Dw9ybCJ74CCSeC2jriDu/QISgrtpZQzYyQAv9BHraQD4KBEvhBHuRh+xoxCxiRFzhBEqGnsMKiBzAilzRi4CCip1ICvVLCVRRkEyMCFf7BHMBkpMwQJXBhDY6v8P7h+bbsH6js8VRiv8SCDynC2zKAsowwnrgPxlqhFXhhH7Zh+7IAGbdBHvhhGyCiACpRQQYLQe7AIdoCGv85Qv4y4hr/4+7+IRQ7IhvHQtEo4hT/zyewoQ6zQxBVQtNoCxAd8R+O4B8K4QgKkRJaAUgUERkLYRt+SxvmYrg4YxHYgBNcwKvGMe5c7iRe4Rs34gvCUTVKESQu4BMvAgAYyCF2ryJSUT6UCgghMB0/Qx4cQh45IhcvYgKPUR6PIAtYkgsooRNaoRN4gR/4YRWYsWtKDivGkFD4ACTcjyIaclVKUSI3YkwmoqwmYhcw8gtY4/ssLe8IBcyiLyxG0iLEICKOABlKciLaICNiy9KQERmPgCzJchuOYAiowBA64c1ochu2YS44wKKYQUUgwpoAqhK/MCUC0qvaSz4yMSX/FOsfIPIr1CAGyeMzuuYFAOANLhIAAAATWIAJnkAGCoAL8iAeuiATaHCpRvIkN8IrIUIMQtMiNK3SVLIsWVIMtoEZDDEmDWze2GAWIIkBnmAHMOENUM8hrAkGIKIieXIjeM1q3MCaqucxO3EsYnCiPgJduqasiOAFMOEL8OAhH5MFZOAJSIQXXuEVDkAE/gEJ7MikrNIhsBIlzNMk5aElj0AM2PMI2uAI+KEer04mzc1NiJEZvDAQAMr//oE3B4USQgu4RMLIQkxL/LIiANMitlE7REYtFqL2OAMBBuAfSPAh8cBjAEACSuAJJnM7X8EBoEDQ0JMj+OEfvNJESfMi/6YvHslyK8VADJAhRo+gGS2hE2IyJinhzWbyJggpEUaQF4KUEhKBwzKCMP+ha4DzIhTUIn5JcL7pHxDSIYqyLBgIQwUAAFRAMj2UIR0gHuJBxyBCPAEOGU5ULMgyItoAGdqAH9RURttTEUHQRm8UR/ERH99sR3NBGClBG4xLSf8UUQBgF/DgSrN0P0qADzoAFOjgFUCBBLbB0ZBgpJSrIt7Lp1RUJOIJI0azTNu0TLFyNM1TEbPQ4vYhA+QhBe7RCqMSUFECAS4sSVv1HzxgI3yyI0giEEAAoFjADX60BXgB5XTUEJqxI0qsPNqqMzAVIuSoTOVIjjKiJedRIpT1H/8gwCuv9R/WNEZDVT7b01sXEQs57wmIlSIoy+2OtCPI1YweyMkqgsg8IgVtTyMl4l29RgAs4BDEgV3+gQ/44PuE0dz4oEwdAgkcglKXik3HgitFszwdYmAd9h9SFALWVFtlVEb5IUbPchv4gfNs4zc7gkIvIqxA1CHgTSxqxSGyx4ww0qdoNSNuhJLcYAAQYALQZUIl4gtAQAB6ADfGJiKCYQpb4c0ORtAe1jPaYDQhYFFBgSImdmLbAGrblB+20ib5wRgC4RLdwFoUCGUpQgY2BiziJm46Ymo4o2sbyWU1AgZggA9koAeKwA3EgQsGYG7/gW6JoAe+YFB34TEFYAT/iPEetctG+9Vfq0AEfERWVWJgHxYZSAAiSAAZnDZyJ5dNkcEmkWEImIckFOljI+IDMCJktaNWzhYielM7+u0fbCxxK2IRDNIgJQIQEFRFdG9t39YY5JZuc5cL8BYEQAAPBtVjLEBLeytI/dVfZRIN4omZKoxax8JoVVSOmJYEVgECqjdyP2kVtiEXmEci5nVVFMghSLczxJAidIqiWlUCCMRBI4LQYJciemA/WCAKvuAOxGEA7hd/B4B3fXcXPEYAdkAFYmHzYqFfAbYVMqdgV1clSPNZIeAKMHdjQeG3kPQOcvMNduGCI0JrRfYfjAFG3mDuFKTfzvdPTwNKKeJd/wFBOCEiff+BBVQAE+5ADuaWhv1Afz3hd/GgY96gBwhJiDzPgFOAPMtCAGXVWSFiFeSBzbhgH7RhG7jAElAmEEiCMQMhFkxXIjyMVRUEZcV3LcjXIlB3YsBYO3rgEsNCAmC4hwdAG1aBC+SNGbhgFtKMF/wgSGPSeFlqLeFoYSHCDCRiTEMCWT3CBi2CUhN4RgZ0WTVCWR33Wf+B3sRhPQyMF2YBWC/Z7DLqQPStejZYgTcibX0IVgQgCojAD8Th5IJUlXOBCnIBJmGSLdeScf7hNC8CkcGkYG8ZLBz3H3h5Ih75JLCVNAcWmHs5jqoXAmoyA0BwTTgvSAnKkxPEi/+Dq6vCAigVxHtRIkdASgUYKBAOQQ7kYABYM0gtYR9qchHBbQj2YSTloRmHePs2QgAZDSwu5mJq0LHomSJymSPyoCKotXHpgA4igmjDAlslopj/4QpIAAIYWnKTmRkYZwgO4Xpi4XPlo99CuDwu+iOcrF3JggWyWXA8WJEU6YQ9AjkdgiXEgQjCGQGgYRssYQiI1XL/IUYdohA09R/WcYhzsYh9alHpwJfBopiNFqEZGqmr9wqQOQPkVhx24A1OuiJg7x80GnYIACIIISQ+GnasGpPEonpYAqvlgADCGQfeUrLK9FNJEiK4zyGMUD3jSafzYCe2hJ/BUyPUtSKKmZf/D0agmdYhhlosgLmhVyGpHbp6t2EJxeGCBVWqIUIBeKiqdwirNaKyJ4Kry8IT/oEaz7g7ZHdVsMAh+M8hxOEDqmAIFFk0y5QrC2EI+PEfyAAHboAMbGAnCkHplsRtYruuHWJ5HWIFmmBsK8KoGzqh/wG4gpoOQCG3y+KwG5oEDpsZt+EQSOIL9E0wKyLPeqiFgmt/JMIvQRslxDhBMlskBAAPAsAXFNIz+A+racMTdiEQqqAfJWIlHQIHmmATmsEZnEF4DLYZ/iET2KFDYMEhBsEMnCC/inuhl7phM2KpjZuXH5mXFxUKBDoP/Bm5LwKwKQJyqxWZkRmpo9uwS/wK/8ThGQRgbw+oIr4zjL8rTC8CtB8sJbgXPLw6NVLCq8vjDDQaBZ7hrH/rWSnAjs5BIpJteAK5PAxcIqjBCQqhnXcaPbGSmEHhCoi2eStixAXbcfNAoFchp0ngryuiw5v2mKv3sBdazCV4CAjgBXxBVQTAF8hbIlyc2NCqQaTjErL7QMw7JXYhCqpZOi47gap62ALhGbAAB3CgZyYiwOmIHph8InS5LCR9IlaAGqQ1WtcTVM00W8VcqCOWIgr6kZ81uk8d1R2XBBx1uYfgGcgByFdBoOkgw/9Bw+Now5d6qa93Yn8LFOYAFEIhFIZADAk9IhAsIsj4kzdCFTAiEswb2f87I9M3ohH8HCToXCx0Srwrorv/AXzxWxiSTUz/wY4GASLsXDUsXSIGoR/OUqdt2j230qaXlQ5WIQ/m4MN/eah9OdUdNbodFeAdV6CvAAfI4MpDAbhEQMOXTIIlmASu/C3FQWaeAQVQoKs4+nNpY3W1mizSoNn/wRsmQoW3/R/YG0a6fWLU6h9SB1YUyxUc/RxgwcDN/R++sx8cYrdRogb+IQlqgB7W4RyMfB16fuctnebPvRnV1UW1MlQPGhTIYBfoOw8M+2CMeiJ4GdX9fdW3HuDtfVHj4R9wwAOowQPEHpE2WzAFAHVWviI4Xi0CpYHc/kAuAe7DJORZRbQ14gz/IOKyV6AZziHA/2EdauDo/4EaqGEQEv8fCl8jmBwWgObnK8DI6ynwHcIfzkEPeh64Fz8iqGFfVuEKcporkRY+1VRNrdUhrDzFdwEFMEAcrgDYHVyhkfhxHVfrAz7gvXy584BWLyzTXXbvK96q/dLawaLuG6kOsiPHI6Jda6GF9v7Y0ypsNyI1lp9VpgcjWkgwnSgTjPwfpCBojr4GDp/xN0Lmk4Ae9KACmiHAK78iKl8P6GEFLJ0acCAMAsHi+zF7R59iAaJNGwgDkRkEte1ZgF2+fAVA8UwcjiurQM0BBSoPBBKrSPz7+G/Ovzx0Vq3ahqMKuV00QOJwCTImiJgf/yPRpEnops5dOnv6/Ak0qNChRIsaPWpUCchA/2qB/HUzDAakRa1RBYriH1OlV7vSvHQzq0tXev5JaSaswr9m/yqEc7WiBsgVIAf9g/VxEKy4K+gJ+/iD7UdnawMTPVehxl5Y1P5h0EEjwJhnFIaYXPUP2ZE2yCB0LujZM6hV4hgGiLwLhRLVgZ49q1JFnMQh24bgEEeAUJU6H2sF+Mgz6Jl/WVEE7+rLqdflzI2eAdESbPPpRK0Va6rzknJaIBFxpa7TGiCr4EGKvZqmufKWTD9O/XjjH12amVzVWCd4rZ51IGus2FtDDcLokd8/59BE2EfN/KAggzSxdU4z5zjjTP8z6zA2CAU6+PKPEmFg8UwYzxCAgwKr5NHRRleEhswVBiFjUh7/OJTaCyjcqMONpinxDBZYTIXFR9/9A5YvQQp1XnlKLolUeyAdN10YPaX30RrlXZfkjBz+o0pPW/DGG3PkgTTmklleBYhPZ97EHVCuuPLXP3qsMMg6FRwYFJ5r4emMnsz1+VEm/9BDgSBN6RBmGLxR8M8NZNzwkgcUXXEFDtuQMYQ4FDyjw28g6fAPqKBq6VQdioYhJW/f1XKJp0HNRFxvTM5KK01t6tRSrR9RWeuWR4Wp63TBjUpVmnH8kyZI3BR1HVBm1EDPICvcGZOfILGV4EfWNsfnXGutgEH/rkMK5Vsk1xUTQLO1+JJrktL1GkkjQ427pKEfGbpmsDoVt6SU+k5nKLH/BmUTdh/lSqs0yULyUzG36sToP2Y8W6CBIKnV04HZWqynxjRtq1OF19YwCD3nyCXqGcAy+891tDil3EeQ/UMDDbXErJMQNDUrFMIgyTtwziCRY2/QRoPHK1FAX6WEJkummexV1vF8cK2p/HR1Ni3LHFOQTZhhnxQWV+vTgRiDRFiCEWqrk9iD/ZSfW9NK8ZcgTtELUsQ90ZINd7R4A9KWLSH8cExc8e2Vr0cP1ZLeiz8e1BprwAESr5RTVbiSJ4DU5U3HxnEsdT7r9N5V0lyDCFHcbS7k/z/UuJLE2dQRhu1NE/qUtk5JhEOPWsKAC/hyfVMNuVELKEm80S2hQ9PVHyl+lfNKTg4HlZRb+Q/2RTmlSufBLg0S88UfJc1H1jAcFC2InIAIDZqYsUImwsTZ1nIg37RxUeusMC1//2SyghO0RGdIQQfimpW67nyEdUwaHVGyAr7maG181/hHKi4Ikqh5hYHlkVxMKHc5oqjiVrRoE/NCxyTvPQ0pmSiaTi4Xh6SlhxunKwoSbhCOJCThHzssD8jyZ7ugJGEQNcDY/MLhtK5obYI6SV0Cu6ckhOFsKBxsTpqmuJwKRo8mULkK+pqjvaGE8ScaTOD4mCMvDRIliT9JT/8Ih1I+aRyrEeoLRw4/Qg8eDuxssgvKOua0AjvFSRiuyAQi3PYRJHQlTaro4hmDEsGgbAEokQwV54iSumRlwxqds0rnjlcdr6DvBJCIwL8aQJRjdQ+KzFHkRzZxNPFVUHpGcV4akhYT7L3RJ+UDSRwiYIP/6e4jwvDfchTpSpr0kSi/S0JaQLI/OJ1AYF4ZYQQy98ieaFGSbKSKKpDQzSbGBB2a/Aj4RAUSUM7qFP/4YjZ3dcmYRKOVRgNEKuIgvo/QsoNE0UUaFkAGdkisG4ISFEgGWRYlqSWZilzmT9ZRTPr9pQaucIxDF5dPWpnyIyjsifyMYsaYcFBQeTQoF8P/9xE1/oN1DNyc93QxFBUKhQcf4UGCNvrOm8DBDv9ghU+qOJ2O5jSXRpmnP8gAEhuYoRuBKs9Fiamkv3QDLvwTGwcJ+I9wvlMVDIOETMuD1aB8NSag1FlYhYIOVWyzJ+78iRlDipQI4DSnoYMpTIFCU6A8VSfHSg8uhyrGKoXxDx9ZKlN9AsuP7PWdK+BdVW8itsgWZZ+zGitQTsHOmgq1OZbtSkZvIteuzlUarNhlPLn0WaPM9Z12SAMr0jBPO5jWghvFoE9Wy7B9coN5zLPlR2YLWKB0Q6Ax+YMizGBSnWRih93YBH8Wq6se9mQTSVCqDicphS8eTy3qHIpPiZLZ/+gx7BSU7Ul4U7ictl5NeldbLUiuFgef4uIf871Jl66mVqr4I7gfKV9pv2venvD0Jw6SHoD/gY6+Hhgp4ADJXcFolDU0ABtgUARNbDGx+fikGxbuRS/AEI7n9oR+QSHxUC46v38s4LC9YMd85CLdo/h2wSBx0D8clNeYNJjBVOHVsXZslAezQnpdvcqy4rCs1N6krTrxKS1huiyaHG8BUuhulaIRjfMOlXKy5TL5gOLTMP9jnv8ARxx0sdmuAHk5d/VgUboBBsJ+hLDGdUIIfsLUFYggGaQgxT96kQx2hEPDMdlhYoUS458II0DO/Icx/7KOcCQDJH6+YyYK2hVWRMC5yRb8AWbDmwqf2tWChaHOfE8RZpj21StCBkmR0cONODhP1iCJAZjHDE+afLe8oL3JNOBQX/6CJBpjbOM/dhqUR6A6s9H4bpq7smo4AJdWPAjmnW3xD1v8Advw+4dcNvyPbtiAHfnw8J/zoRMbdGMUB1U0UOhHXVe8jj9l+UsmzDDpf6D7z5NegQ4TfRUa/+PBQDmza5nU2n/ANiZ/Zc7VtPwP98rztTQ5+D9QyGuFz/MR/5iGg9MzT58COyj+CAgAIfkEBQoA/wAsAAAAAPQBGQFACP8A/wkcSLCgwYMIEyo0mO1gvYUQI0qcSLGixYsYM2rcyLGjx4kDPoocSbIign8TNjYoWZAby5cF8cD89+Ufn5kbVUj4J+ESrpdAcBJkIVQjFwb/uBTluHLpzKbHJjndWFOgtzQHAUzdylWgqjGBlAhUoWLHlHLVAFSbBGBSWkyYduywYCHKv2e5joaauJMloq4cGSB1ascb4MMX1yCWqPhfAIiNFyNW8G9VyILKBlYT6GWg1M8DO5f08mAEHz4jDqbsCOOfDMkwWVS12HSjvY8bTBF8BbvkSsWNuXnqTZxkKD8slv1TPjDzQq1S/7XFtLDcsY/X/yljDqBcrNXFwxf/9IVV/EQOCduZVxi5oACB7RUWKPDR2mLK/xLkP7iy9uFy/7DgXEFsAaCVQJh4UY6CzFFk3UDLLCjQgsqQVhCAmw20gx//uLDRa+uFKOKICt1D4okVPTCQigXFkgswhgQzhUADkgTgPw+U06BENRoESCOXYMFJeKL4IAqKSJ4IokKpuPePifL908FIuiQJEXj/wDFQLDwK9IAKfFSB2j83/jPjQSxCSKOXmbUZEYAATpHjRGci9AY5Vuap51ZE7EnQN+LFx5gSxlhUWiyBJFRmmQYFReYUIxgywlkQlfPAWZFaQsUIl5Yjp0BT8BFLnQSpmCZBAOxSnp+stgqRBa7G//pPCUvIQMlALQi0Ggp4jjVFCSyQqlAOI8CZUJpTBIOGQCOgUcU/VaABTC5kFnRppCO88UYwhhgiEBpUDCFJE5I8s+w/3HZCBRVHfDJEMNWWumJoI6gg3T8CaBtMIIJuNU09/SaJn6wVwSpSdgQvVYJATFDrBx9qGJRaQSPkosKM9kaM0MJm/uOIx1NM8WwTVZT8DxUCSXKLQCs38c8t+3YaahADUVEFFcAo0sTKAvXRxy1NDIFyFQaIS9AtZADz7AjBpJABjIZEDOk/o3L7zwhVPIPOQCtpieQi/7DxDzNYwKaffhJ98IFAUybsNqvoDcSFUv9YQu0/aogjEDi3PP+DdzCd/DODQBrj/Y+9EDHyzxAFYWMHLo9XWQUBVVBwyy0+dxPCAjHYEYPLB+FwkBMCKSFJyuwMMQQw6wax78RDj5DaCIGMQA4FEejJQdxvH7TLUqX0DlMkjh1EyFaelHEQ3QJlwMu0lHRiAC8GFBRCCOQagfLJVNB89Yw5QEoIzwex8g8PktnSBBh6CxREEChnIBAwaBQ7gjG/rHHbQA3liZTXbovEe6biAIGMQ3gYWcMaAGGlWQxGILPgAgtmkJpbVaQQAmnCGMYAupc9o2/k+MU/ftIRQAkEfRExHyvMNxBJFG11BsjA0xIyAjVMIRbPYEUDGkMLgeQAIxzYBgL/hzgSrz2EiAYpwkAMdhA7TORII5nFPlBzvyCkABgJwSJBvLcQEspKUjOKBTnW0ABE9ACJaDQP7xC4AxHtjhNcyMUIBvePW1Ghev8AFx4PosU0DsQS9XNECXIRizKAKAdL+OFFTnAYMj7Cjy8JHkdOUpELEOSMEqHPP0CwEaScYiBHjAjiHEUYENxkIYTAAhZuwAcWjIBjhkjBQGQpEFoWRBLisAEFKOCOTCRhBVv4RyZgIRAbdEQI/yAdNf4RDlesYBAUcIUNGDeQPrKEZq6b0QUooYbwQdKPWjFMbDJiyScgUCYSOQBJ/BCFZ4hjBiWYWC4MYEuFkGELwvhHDb5p/xAtVoF2UzCGMXyhwH/IoSAP5OdA8jAQM4gIYThBj9gEMqSNtHEpivGPSCxESpxsoCCB+MA742kTS6RgCAbIAkJicL5/sFShCsEi/P5hCDRIKhA7ME0LJpCLVJioh//g0D/mgB+0AcacME1qR7aWkDMKtTfKUwgn/5GoQjgBmW9jIWxQxlXuvc8AmqopH4DBhTw4QAMC4cKtREgcC1xUJJxkoqyI8o8XHM6PexgIXZWaMGoOxK84keUQUkDYwRqWsJbohKhG8IRchAEOAeuID3zAVyU6xUOH6YJH8ooRBh5ENCFyRnEWgJAVwER+AgHsQhhHTVvWMyGold8QZEhbGf86jbCdCMYMZkAJcYhjogQBGyR2OBCs/E4gd1uKBijLkQOVxK6Iu0hHKQK2gsh1RK3h61L60A1bfOIf3wWvDf6gCHaAVyBG+IcRSEGKXoTXKSoViDwg8tqC7BEhWchAITKQ3/7Sdh/oyiMXtMEMNrBBG9pQCuXEUQVx5CIXLCjB4GbQAl5YMk94qAk6xbPh3r11JKIZ0GM0YsGuvNQj2MCFP74RDjCk9x+2wIZAHimQd/jjke/4B417F98sHMHHWQhyIYLs438YwBCt6ASALWGJ6RF2HxnYxxD4sY9E5KLESbrodXvj3IVU9yLJ3cohpuKIHRVkLzN5w0HCbJ4dG0T/xhghw0LiK4Z/1Fkg/DDIEWDShoG04QhiALSgA/1jMWQAkGhQMiUS1cZEHaQSqJCkQNQ5EDUvhBNr1O5EKvoPIWr6ak4KDx1kMZBM/AMJp/60QvoskiN4+iB1RkYbZC2GNtS61kdAhhj4kYHqITkXfMhFK3KxTUq0oAXbYMYqtLHsVXCCE0MQByV4wYseZEjVEFkVtjWC2X+YgyA3IAkedoEHPAgAABZgAQv4IINEKEAUDoD3OESRDAyMYQFj2PZCSFASCPgbAvyOSJ/bMGtb6/rgR+DHEY4gj4VfYRXxSMcrCOARTqeRePrGyF41Et3sLgQEKKCJTAJhjFjwIRG8/9iHFClBiSQPe6wQyHjMC0ICUNAhH04hgc7pQId5gAIUq9B5HkBBgm1sg8F2oZobJjCHpobIrmc4DCS2jcmPcOkfW84IrL7QZYH4wQ8H9YQxiOBgQhKAFxngwj54AWxDdMKkzNAzzjfRFdFOBAmkhQjdBcIIZPxj5gkJOMABfhBQ/MPweaADFOjA0MYLhd+r+PviLMGL3qZc2atg6CvyoNmCHPcfnyfJAElEccQMJ+mX6I2lk85hAMhkgBQQSLhLfwYU2J4GvkABAYawCn74/R/8MIMmKjAQu/+D+BU4B/H/sQ7A7HMgph3EP1yxzIGIYb4D+f0/Zq3rgf++DTqvQv8hGH+FmUc+8AMhOtHzQAL2E6QXA+H54hfveL4HnOaVYajhBaJzouv8/zq3CquwDYVgdNsgAv+AgBHhCxahDkiCAQIBgQgRbv8ggRYhDdeQepcwYv+ATtfwDxhHEBxYHEA1EB2WJGtjEDSQerUQeuA2fcLQDOdwfP8gDMREENXHEaYlEDWQT/8wgwZhWjd4ECJwBZ22CsgggL33D7lWEKzWBhAAhf9GAoN3eHQgDkoQCGfwAmcQCO4kgPHAc/t3EPy2f0OXB3kQD2qoAKFAOhQoEFE3ECH4D8UwEM8iEKVHCEowehlHEmkgDR0RBwmBTPmWbwaBCH8xEGFAEo1Qh43/IBCPKB5VchCeFRGqIEIMCBE3cAMrIAUDUQNmsAL0YBAVoAf5RA87SA960Az/4AwzCIQEwYqsOBHGVxArUAM7aBCqpDc4IEQ8JxACOHhUOIwAp3MQwAjGyH6MkIZDQAM6sIgQiAVhsIgDkXoH4VACIToEEXIUIY3/MBwwgVWSUQv/QI4KkYm9AhhQsgba9g/tiBFsJRkfuBBiIRZbIYgfEQKu8A8r4IMV4Y8HIVrLVxGwKBADWYMGIQgl+A+aEBHUWAvkWIfmmHqkpQMFQQO1QAMHIQhxSId70kMRSRyJiBMAqScWeSK0AAgL+RFOJBDREBGTCIj/oAqqMH3hkAQC/9ENBNF8CFmSFLF3B6EHBdF8B4mQO2mQ+bSPBuEKnniSBrEFppYJwSQR8XgYlfgPgMBIAmGRWnkC/cNUCDGVCdFDK4kQufMPWyCWFpgRyIRqEDF1fvSOGEFabikRqaAKcdAkFCGTeskRblmLHAEcdKcIBKEIhJkJzzcQOmlq3eCTgCEMOGmUB7EOthCKmlADrlADcEmDF8FSfbkQVVmTFhEDU/dJ4EAcWvkPnrgRLjEQnzkQZ/kPsckR+ZRPRRkRL6mOG/EIuYkQ/jAQKYYQrICP/zANG4EVLhEHrCANP/FJS4ENZmBMIVAQNuBQOpmTCHGd/2BMApEPUJAPvRCeA/+RDDYAlAgRDv2IEek5EEngCggIf8mAc1DADmbgTKW2Aq4gDD/wSZuZbQLRkgahVV7UG7ogl/8wixIBoObjnAaRO7kji//wAy45oAQhDZP4D6dAoQdBQgBUEc0goSPSAP3Th7KiSCTKEgl1EB05EFpwov+QohoRWSxhVyRhnOL2EvbgDZb1EZRBGUZlESbigsU1ggKhbb1ZEUGxJB6xBk45EEswEAIgEwaKGEhhjy76ESPKHhnhDeKEE43Bh1q6JqqWCFSDOBLCGRPSEZuxIDeCOLHwpF3BMbFyYR5hH7ChGwIBDVe6pweRAKvABmsDWhghqGIqEMeQIQiTqBSxGdX/oAxX9w9kGjYeoaR8yhXApRuowBEWtx7BAY4C4QaVChE5IAMtEF0jcW1pOiEQdRGEKhARIhDRAQA9cBJssKmfhlShChtQgiSa5BEmMBWfMicFoRxeMCAowwLlYCkKwSgWoRYL8XkGYiCYYCD4ci8A8B4CIAA9wDwUIJO5+q3Cs6uu0gF1IBA2ahGQYjeG4GgHASCnYhHK8K7awawRUSP0KiJo9TZo9g+Z2ioOOBK9KhHvcZUI0QG9CqoTAQd2ahAXShFP1RtTIlS5MhA1GV09QkPeYibyyiPVsAsA4BxBsbEHISck6ykGIbILCK44wWZ9GInw8RILWxy/OhGpORBY/1Y2ZSMQ7AoqlaIC9XKvA/Ku5TBHnDIFgcAt3WIIO5Cs8YIjU6AGsaAGyQop3uItd4QykNIKZjIDnYAGTaa1x0Ip/7AW/0BQAwFAJrQRmQYTwEUS6vGtT5p1KqsRFlkGlUAJswNqI+BKsoM30WUaE0MQ0+UlU9CiKjIjpiInsVAFMgIvBFEyBkAGxqQIhUK45RAIM5CxBOEsfdQE6iM0eURTODMELjOdBBEyI8ALlhC4KyI71XBRz0AOJ5YnurG2sDEwCqE2bLMncpqJJQGg4IoUXFBhg6MGqZExAxEDz4BJkUJHBTEjzvteCQEFBmEDEIhvxjC0NwEuVSAJQ6AIK//TByEQDoogCX+wnYpQCBikOASRDP/QBHbwC00ADFg0BEdATesyAyEDOJ2QuUrzC3bQFBo1tzgxVQT8EkTqGgIxZsQxAUqxD5RAQSPQCpZgEKbLLX2EBolCKvfzC2mLENz5DwvwSJAzQiZ8PjzAA8DLA7iAQhWRwu4wEE3QBIVwOt1jU/8QBMDQawQxBOQADh16D3N4IuhBSQcsEu1xpN+0or0xC8hhOMFgANgUEfR7Uv8gCWQgCalBteFriAuhC1p1EJOIC5PowheBPYpwBacTBFKcAbLUVegyBSrQA2EADvfQFGugChYwuJcmGdS4px73Eh2KEVF1xAKBpy8qRRL/bAxYNhFchBBgnMKHUSUNawDhIg8ztBA0IyNURQi/0ACgTAsqYKL/YAWG/BE7SjC/kRGUChjvQR0X2xu7wwFswAtRGwwVbBD3pWmWEAyT8g/GMAbZ0AOFTDB06idgmie2KxENeyJ8PBMfrBDoMQu84EqtYABa2wn1JRF9VD3W1BFVEsb/EHsSscvl/A9YlM45nEeTwgcsVwZlAE+s4jcBmwu4esoUwQC2SjB9QRKUFhGPihCYBjZVYMuvNGFNZhCqJRDiIAWn8A5CSRCjOBLCMNEHMQjayEcz8T77MiuU0AMCAJb4nEYwShF3IwDmuBEFxBHHXBEPcQ8EuxVyEAUg/1AFlhALuyU4JlU0f3UQ2zCdQzhE5qwQKOPL1TAFVfcPx6NUb3uiYvNlJDKPSzEbU1HTBg0vhWCPCzCbRLTNEuHVBREEaDDWY/06FZMIh8AJ6nQA1HsQbfMSlXAR0TDIHWHAIjIYH0UR0EUwVK0QZ3QHA2FXQqoQk5DM6xGbXI0RiU0S/QkRC704RUFPRUNPTmPJM6BbhtBbQlAl4goTzBURDOw2RWDYJIHIGNHKGAEPIxHXFUGcaGoengiYi/0RDhqhFWFaGgoRGCQSqkVNqKURs3VbbuzGg2UAfLBbuSAOWIVCsz0QNGY+dxOpOPHPI80RmtV5GiGnI4GyHKHdHv/R3FPxXZ9ACp/wYqclGfklQ+nNX7Z1aLsVDLygDZywAWzwUfRNBKrQANGQmmbxD3twZcfWAsv8Ecz12RpBHQJxIAjuETTaFUUAK3KrekvRqkr1m4/QDdKbd/5gY4+ADdgwBiGgCDawDt/wmyESXwQB1gMRZP+QBUMWZD+WX/uVXylwLinAC7qlW8d93BImYRQUC5QAwSyLIgaTYX1tHm30VtVlClCdSf+Q1EuRIajKElOeEE2HGHVZHD+RYwJh4g1VEYyTBdiXEXXGaiSxZwu3cEC2Zy2+DYcWbJbAD0aXAdsgD6uQAQEtEmIzJG1rEE3tERG+JJnRda3C2vls2hz/ga3/sOBpNOQCkeV+tHDrYWsGJwaWHmh/JgbMsA/dwgeGwAe80AK5gFN1cgGV0AFX/g+fPQwa8g+WVhHUvW3MkxTguq/i9gblNhCt8QQywAtzAG+iEA9tvQCQXhCiJVrgfcoEZ+YEYea0xoR2Fu1Rprqd0AmtgGSf3gqefu2t0Aq9NQIfVt0ewY3Cw+gcgbAQ8QYokOtYp24lUAKHoA2vMO+v0AV5sApXcFUCIY7bFnC/yL4aweYIMYwkkA9EZ4QE4W9QuOyUXmu+xw95kACvEA//sNL/8Aq4i22C8A/lqmmWxroWoWavLhB5vk7/MAAhgfIDMNMvYHu78Aap8gaM/7x2vNAJ0YNk1m5TJ8W+XgwbgHkQ5ukUoOBzimN4YziGFAF4BaH0/EYCyLANXMAMzMAFhmAMciHzJlcAQ2LrXPEGgy3uSFK5A7GzMCEH4nAGILADvpUIQc4MeZZn/zBfYy4Qr1YIV2CEYpkwyAABPHd/9zfw/Pd/hzf4BWFzisd4/zB0SM8RTf8PxkiMqwABSMhr+8BkvLAKqW4QvnuiUh0RJxgRXVgcGDfy5jF6HLjU4ywQ5Pw71ujqmwSHFIcDW1CLt2kQxX4RQV0QuT8Qub9MHpB924cQfSZrCy95jv8PdLANY+ALgUABIgAK9w7wAE8QRp9+JNALPwcK2P9ziv8P/dBPByKQNZ5AAeLQiw9HdFYICq9AB2E4DzxHB+lAflcQbc8wBp/XA4XSbXtaeqkGEP8EDuT2r+BAhAgjJUSY5hrDf7sEooBYEUtFjBkTFvsHqGMjjSE16vhHUeTJhAsy1qJx8ga1Gnr+VaggrIIeKf8GCXQVEpbAFQJrJKmQ8IezH+d+oNRTA6Eralv+tQyEhRCFKtvm5OEHQSCygW3+QfBKAoJZtGdXkVhFZ86NM+R0+KJ7hsLVqx/uYkHhK4BAX5eqDPTwrzBKxAhrJXxxMfFjyJExvpBc2XJIkpc1a8wmefHmxDRUVqZAAeM5kUUFOvvHGjREev+CPhb3D4v/X7//AhT7y7FYS4FC/gUC7ithGISXNtda+PoycufRJUvJbLnBwHsD4SSMhhjRiYG/VAmMId28cOFTzYfsniryFjMrksROclJ16n/rohddYTO/bCQGUuKkOjbKqDqBEFkPMeEQfI2jBRGjhZbx/oFEIHAinCmxNUTqUEONpJBJk3/SeywOgXTJKJVTTmGoQgYREiax7Srq7h9p7PhHxRhsYEQRRWz4JxOE6usGtE32EyiJ+v6ZcUlhepJNIxNFigDEgS4M7x9VDgoJvIE8egiiJiFyD6UrK3uos3/ArCgOGEWKMzIeBDqlTixRkkZFgXS8LM2B8BQIRVbWQ5FPy9LA/+hDhKZZY40GNnFCkYSAdGK2f7rBVCiEevmHHVvW6UaY+pIU6EnpMhmEGvlQfTITTZ0YKB9ZBVLVFdcSakYkRBkq9Mx/XMwzo4NQRPEyRJfSMiFnchJIpQqcTcjLhLRclqFo7IgGlxsTcg/YipwJcFjJGvDIPAHIVXdddtt117LaBOLiXXrrpZeyy+wRqDl7XytAIBn6TUgCPEK6jt56GJIAo3RxFHggBDIqQTIiFsTlYYYWkc6a6BYWqAiMAMBYOSA0OxghCDGuiOAIS15wYpUhmvefiJVgNGacJeM3Z4y6RQjkge7geWiNWBjhnxFYsAAFGgJRIZAdAnljl2x02f+uw3BESCiBgf5KyAqMBsBSUYEeEUjsdxkgd5qdiY5QmUUja7uRk93u9wKBElnXDYQmEbkaL8qBqJpJBKoGocAF8gLwHVRg4YN/mBnuH0yWwLJGgWAeembEmCgjMmDhAMludju8ObGGRY5wGkW9Nph0iCqOjoWSF//n8IFw/6fw2wcSXKDf/ynHi4yUIX4gTBAa4Yl/NBeog4xQ+ScUySyH/aRWLPtGII4h01e6Da4Xf/zoVtFmPcD/OR4h3RETvBw1mO8gl0MKOEQ650VSm/zx2UgImi5oxgV2GxD/cma9gfhvB5ZJ3vAwcoz2vYZ4XmAB86KTPwPa6x3/qNtm/Af/msNgDBCmS4gnMhgzKyyMDVwgBNw0g4nF8S4jwUvM+v7xAOFVZAe8EAgnTni5HzKkHRnkV7rO9b2K8E0gCNTIweBwrofhYCBco9hAoIcYG2rmGP84hvEE58IcRiZ4NBRJIPwQPstgUCOcC2Ib22g2jPxLIHdQAWQ+IxDX0WsOGTnZhwomELxJB4w3nMIIcjEDBw6ucABQnRe8GMaMbHESw4MhFweyRYFsMXDrm2DyEsILH4bwJEwYSMAiQwg3ppJ/SFSlwHD4gOC5EIeO/McUZvAPSlhiBlM43iA3Q8t/LOMkABAAMQfSHDYNKg5xIEfE/nGDh2nAPKdrZTVzlh1V/9YoGwAwBkNwqBFDWIIKxghEOZTxTengUJjr++YDhHkSMrpNFOPYjDMxJj1r5lOflnFhLHJhiGAkxJeQFAgsEYJOyeDQl3Cbwj8G+bv3VeRaqeTAw/BpwD1S8TWmREzDNCJHgJ3kOtvDSAcz2IEWJIQcLMghQjMSCD4g7YYJPSfcbOpQlDS0HC7dZ099+hqPIkaJiPkCROJgUsxlRA7OCaB0gIMSF46gFUeryEAhooxyYOJw5RhBLFDygCnAcgqxuOVBfRfPivBOZLSg5k8F1la3xhVnF+oBZJKmhoFYdSDfhNtOhXfOQgaDD4bAK0HBCtZaAk8NZaWCJYIxBciWYP8K5ZhCQAEqvHi+MiEAAEGGEnIyP8l1WCRsIwj+YYGImGd00/hHhxIm2pPkbwIDQVtLjFFHgeC2oVUdyAioipFBgnUEhjhaZf9hiH8MBiI4LCQfRgCANwz3H2gQCBokMQQqNBe50qXCP1IADJF8cxKBCAQKfmEcuvxjDIJSlyxUNkTLKKAi1zEpbE9yiXOxFq72TUhLmMC8RHChBQL+x4D9II4oCISszv3HDHCrkcmGlaB5nYIKRlAOFQQDuQipgnUl0d3dDgSyGiYudTeMBioYoBBkUAQYhpBchKDBAENowi3I0F1HiDgWnbiwQ0tmvBGo4HBvWOA/yOHZdiVgUyH/sad0pLgZ+TKEvq0EWsr4y67tsOBzF6AEHywcEjWoYAbOc9k/tGDmf5QMCFMos0LDOtYqBCOgnRhIFYAxBEkMpA9NOOiINzwQNNhZEZK4hUAkAQYwFKK7AjEEnv9xixDcwgbgFYhxM0CFx1YaeL8diCo6dDDlbI5nUUYJR8k3MZa+xpMQqe+VQ8IFXuQiyAN5sEAs8Q8KULWQZWUIV+ss50AEg9L/GIIBJEEGPkOk0CGowgggOwU0IBfFKJaEImr8jxD0oQ9jWMACQnDdO+O50Nj+Rx/+keeBGODSxyVuLUfQCeK24rKuthu1eMbSUK8nYa0+iQlczYVZUILXDCFE/x2nYIhO3LKwDKlCE8jAkFVoxAkh4ME37PCLZwQbxVQYgrjLHYJubGI0DGGEQEqekD/8QhLgTcE/SJCF7lKBCs6eQi4oIXM0RC0QYwCHHQ72Wno/DEWq+4epg44zkNZrf/KaRUxjqgbfiqMQ/0DyWOksYobU8RcJ2cZAwFIRPuECFzyIQQzgwAN3hGAU69WFinTBXpToYgxk+IMt/mFtMHyYCkEIxgjQEAQqpKDlAzGEISShhF617eiLR8jn7Kt4ezl+ILP9BwMs79gZGCLFBjCAOPYxhK8LhM9//oclKMGQKUigCoGACC5Ci5Fe7Sghry9UYnjgDGdQKgR8BgZ4F//9D2AMPgVouLAxzmCHNWTnYN0DgiPAhpgPkmvp1VxIUAUmgzJI3r5QnG+ehGZBeVVUIAyYhTh+G4tbG4DS6IYIeDlvAEsQViBqCEQVnjGGy1xMRWK/TLdCYAtbGLQgSLcMyIIgoDQewzBjUAI4uI4PQYd/yDHEMIUBij6R8AGBwMDKmL5qsr4FcS+EKIXI2C+iYSOGIEG3mYV/4AJeMwQDQIgB1AhJuK4quIU+CIFza7YpqIIx+IUMuZjWEwggDAkeeLt/gDuNqJNeYYRCeLF/SLEswC4D+L3pUoMpUANCQIEG2MLWSibIsEDGgx1RCMOBQMF/KAK96pdZ2IcZOJr/GTg9gRg2GHxCgXjBJzyCKzC32YuBMaAAd4iB14uM2hPCyug9YhuCDMgAYJhCiAgCvnO2rrKZe7gOWviH5xOIMzsJNliEriPDzQAa0lkDQaAZT1QX8tsHPrglYxhAOUyIAXzFf4hBO4QIHigUW2QXJBSIAYw5XcQIwJs5yJqBZ0iFBliDWki1UqyXS2wjM0wIVtgZo2uXZUhDgWGDQxgBNQiohJjFoAM8NFADvMoFHVgDWqirJVpGAwKpXCCdY0klyjvBIAJFjKkoThCHWBiBYIBFKkSJGByITmwlNICsEcjCHsi+f9A+8vGEC5CjdUxGDTEFh9QMrwoJTuACWcu8/3/InqtLjH5spWGjNMJarBZoBYNkojYCv4hclysJpH9gAo/BiKF6DQwYRJEoGDVLs3UBAVISiVngAqOJBR7KvFkcvIrgvH94wd4zRPACBvZ7OM1AsitACKUciFaMjH7syNILAt8qsD3gAzVKyRMaQ1EQwX8wrXzTEHNEjKR7joQAOob5BxWoo5fUCJdByMiwA9MSiQKhgFy4xxmwnBmwBG4UCKIEPuA7PG55hx+QCYYgkstIBnZwhRpwCoTQAz2gB1fAgaU8SsMczM0YNuJrKErIhSVYIO4DS5/6StRklyj4gGZrw39gAcE8CXEYF3VhTIGIjX+IF88EEUuwBGf7B/9jiAUUWAOSWs2UTBi3rIikepedHMGBKLM8gUg/iIIXEAceG4FbagVLED6MEAccCArcVKVZ7M2EAK8B1MYReAYl0AFyQAhPgI56ISmaBJED0KcQgwyI/If9rIgxybrXcIDIaAA3CanxqU4Q6AFeoAQWuKUZaIUUeMHBHDwS0BpqMAN10YSlGBoqmLYZKLJcuKKKqCsHkKZ32YMgyoEc+AeT5JlN/AcwpLdlcARHKCp1eYEesIROIKsGa7Q84K/C1IzuQgM5o7lYiAVyyAZfWKB4kS/qUZe1RM422qMwtIAoOIRDIIArGAXn2CB6wQUuXZAgFYlpCwI0INJgmAFgkAf/OoiHf5iHhJiFSgCROU2MO3qM+4SIvCyylJLSYVk1fbqfxIiAXMQZf4iZveuuIHg/A4hQYAiGI6UEXtCGWUgpCGQlVcrLyYuZdzwJZIwrFP2HHvjUk/CoSZgED7SM54wOlbgSQAmiGRsIJyQ2kZhVwowMwUuBIcjVXU2BXOi7GZiBXCCEBWjGy8BADfwpeXSOBKsIH/oHjbGXV7iMOoWM/zweGRKYXEGIV30NQOlWd7FVyMgAWX0MXc3VDDjXdM0AXrAEsuqqQ6gCdLiOCJAKXBMJbGrIkEhWZcWSZ/2HfxWJaqWcE2pHnrHNf5CW1gBXbx0fcUWIhw0J4SNXgVjX/xTIAES82IvlhYQLVj8ghDEYAOoJWIywB3DxU1XiGo1CjAWKxsvwAuLJVpXZVnUhhYTwFIGwWSMglyxgl0QswJ/92XMNghkgqxaQHBj9hwFyAQ64AUiAA3TYBRQwCXXJU6JxGdSKDHQcmmnVDJd9mDkd2M1o1X4xgk8YCFL4BJu1lyyg2NfoWbgF2rZt26DlBT4QrH3QBjZggw3YWw4ggGuAlH+oBRCYgh54ghbghZHkA17YBzT6BxOF3Ojg18ooAtP6Ixu1DOlUl2fNWpTtqWnokYH4hD/ABmx4hG/Ahm4IBycAg09QBCNQhE/oBmxwo54dCLnNXbpNge5qBUrYh/915IOYMoZgLd5gLYExk6oW6NPrsVEbTR7V/NxPuh2iixDiwSTniN7XiAFniAGGjYx3eARsyD1KEQiK+4fa/Yd3OF1sCF/xzZOpI5cMKIQsqF/7vd8MkIf8NQA0yDxesNtWmIE0DVbBCqcUkFQeCiTmXRAMdFPNeIOByFzpRYzqdcjyII/LONT0fV/9YA1sGEKEMBuzSV8N+Ud1OYJ/OAJ5OIIsYOH6FYie3Qa+4wNLYAZ+yIBtwGEcHgJ+2IbV+weWvIz+DInIBQ1NhYi5pBcILjKBWASSJRrP1ZB1eieMIDXEiKnXQFh7AeHLODmIiN+EEIOB4IcTFmMxOIIzVmH/FGbhIziCSzME7tyGVcjhXGC9KI6ORWCDJ66XCj4hfZ1AoBIICP4HLH4XfLmMpfooFQyRd/HSgTjUBWljiBBjsVAXSkZjTG7jNN4GZuAFQxDgXNiHRGCpIrOAmKyIUqDczdCaI17NIG6XVH2NWmOXQw6JMRyIkRMtMhZjjSBjLOGHNvi6NhCDNjiCYj7jNuCHGzYAeJO3YOiE322BfeChSqiEREiHf7hlUdjmYVgFY4iaKDCGQU6MW/6HUoi4o9sfE1w8aryo6MCDPxoIGBAIC3KALogHaRoNlcjlCdYIFE5hiKjkfxALgv4HZEjmYUYGTBYDedgHYKACQ8iFVugE/99thScYrFbIaDjO6ACOBUmdAiZOydHBiJlZZzLMowECkV0QADwoJgsogRLgAyYgAgWwZ1HognFwU352SK9YDwgo6NCrCF8uaIAWA4ZmYf3dh59lBhzeBjp4sWoYZ8toqrhapgihWp9K6QjZBXh2aRZgAZg+BADqAgdwAFHIAygQgUxAAvzTYsYjAVAQCBLQDIEOC7I4i3wABRK4AhII6oH+6TYI7IMWA2QgbMMubIUmAToYBgdOAMghw0TOCEAgm34G1IqQnYx4yVrGiKn9BwhumK9mgUPghFVYhXRYBYtshVwQATKokqCb64QggbyGCNh+jbKQbTrY676+a7IYbP9k6Iq2WItt2IYEcOBsltKG+Ys86ucI8QM/GIAB4ILoHgA5sM6pxYM3gK5cmIVckOiLzsiNlrdWQANg8OKHoVl6ge18oIO4xoi5rm2GAAu/1gizYARQYO8rAAapkZo36O83eAa+eYJ5UQAqndYf1Wrm7ilSRYmiiueEWHDLqCuJ4KEBeG45oG4Ee4Gp3QUQYKQ3GFUWiAVxYIZtkGh5C+UVloeQuA8QYQ1AUViBKAq3tm2zGAj4Foj7zuuSi+sfbe8IiTgxSAFxsAQu2IeuEwd9VYAfXdlhcXB6kwjSGee0RAwoZwgWEJr1eAECQAg56HIiiIJAOIQhOAReIHOby4X/37xYFUfh2xUINsdldlky5/hRCGAEr+hpjCiLsSABPne5hODxPJgHOqCDfzDv17hxlzsLCFgFfpCH/82lRKAESbUEcRBZKh2IdDEOAcDqBL+ehRidhQAa1hsaKJcIQa2YG6iYMwABVo+CjkuBrpPkfwDj3RyITUACm9iEMMUZaii5H82IqIzvREcGUACFYEcMvebzuPbxPGjvPEBrOpjt6OBzPld0s1iFRUcGZEBErUAIKx4I40hGkBhp+zpkJycaAjCNgVCOS9iFNzCGrPDlfpCKZkBvhNgJLPkJjcD3f3AFDzh2YS/sfyDmgyZqg4brKtgFSZgDOsB2gUBnhKjt/2X/B73W6zyA62Vv72KP67m+bzoQ9Hkodht3b2q/eD5nhGpHeVDQhm0QhyroAWOomCt4UvMQJVfrHiengXPhmDsdiGYViM1uF+WAZ4Fo5fF5qoo4gy3/BzN4EtT4h2Y4h/GMDH4PCcrUj5MYhH4A+H8OC4T4up8O+zbA87OgA3EYAxRQgigAT4on9D3HiF//h4tvdroHhYvvhTyIh3jIAxzIuEB4gUBg9QAIgEggfN2gi2fYTXFYKiJYet0oGDxwHSjvppCo8n5eA2l4CG9YboGQhoGoRIQwDspwkAV5bI2oBW8gnzqQz4TIt1oId4jAARzgd2eQiaCABaeghqqHjP/JpAdhOAelWI1deQxqEIFtIAO/r4KsmIOIQ2z59jreJgVrV3SBeIVtwIBAOAPtR4Fd6H5PkP1VYHhQeAU6IH84pfg8WIU8SID0/4daEQhq+AcTystdaIm2aRvIeWzWh4gzAIh/AgcSLGjwIMKEChcybOjwIUJuECcaVIIQEUEsFB9m+weoUbGNIkWGHPnPF0NX1CgIO3fO2cB1g8y4olejxooVgwb940kQVg169CqcEwiT4I+jDV/+g9lMWJJ/rnwWxIClCgYcCV6tgkDwykAIJCCQHWuWhNlVefKsohAoAMp/YbBgsTpw179LA31RwGEyocZ/gf8SLuywVsIXgfD/GG5sksY/FALHLNzieGJIdHEESluI+DJBQAJFiyYI2TCFG66QJBm0okLTpf+aCaxwVOlGmLgJhhuI4STCG2QGkiFTaNuqK6vUMs/DiG2eBIyUb8MhjoASXwEyCh5YZ6PFg5FCWgMNkfLAweYb0sB48Mz6+PLnHyz9zw79/A3DUfuXiSBsCQX4zzoIDWjSbgTpodB3Bt0g1UCQoTRhMb4UQ8tAC/wzBgroXUZBQhhmY59COugnUB11WATiiQKp0mJhaxAUTWOpwNhYe5+ZZOJDaRgUAUR6rfDPCv+BdqB5URWGIUGIYegeQqfd2GJIJU1JkCpP/gPJi+bxqF8DDkHy/9cJVx6EhGOCmCfRPzYK9Ms/ZoTTDUGb6IekQAUqpKdAUSn5D5osoimQEAVZ9ttEUA6ECJP5keZReQYtoIOJjTZk2WWITkRLlwRpgiWoZi5Uzz8yKmTqfFKIypCl+k1DESDZYOBEQXQamSdhfBLEJ68U5YRkEjTdalKnrd6oin2AoCNQmWUitKxC9PyD6UEdCWTtQp+SqepAhQ6E7arhDrQZZyYNatAPBnXpJkG6KBQNKwMBORK38tG4Rgj/KPKHQGYYRKdBwsiH51/CrOAKka4UOm/ADnUZA0TGQgRxmxSLa941LgqUMUIMLwQknG0mJPA/3iJ0yj8oE8TuqvHG+/8PHI7RJlC6B5FLEH4K2UEjQZ2BM65ALJ8Y8xp22ACGQPz+84cZZqyQxJAEAfxPOCKw09tAwhAsXw1m1ECyQuz804u/mWTiSiYoD6hqvQv97BDEY1o8ktCivu2xQwHWPZBEEm02pkAexxAvjZ0lxINA7kL7D5JtH4SLQC+zcgrPp5Z6uWH3FBTzSDkXNCYPHrOCOORubmb4SJzrwuY/urzsLuojoarQN+GwY4tAuPfr9J/DEsROPgblkwwj7Dhhgw3/5NuNnQglIYyuDRk8CDVRF7TJCrT+k08v/yTDTk4C0UOBKwLj3ZC7KZ/cJuIXF8b6P6y42z6Q/izUjLM1EyT/kY8FnXJKuvRnEMi5r4AGPCACE6jABTKwgQ58IAQjKMEWDUAgXKjgBDPoEBLpBwgbbAgIGriIjeTAJApYCBEyOEINToRHCMAgC0eSiwbOjj4SUIEEBvKFjXAjEjE0iJtkoEAtDMSDhsFDEQyyDMKEySCV+2EEHxEfUUARIj3IoRGrWJhO/cMNCCSiFnPoQAYQBIZaFBcCJliEFxiEMWeM2BeM+IQMbscgNUSIClwlQTLa8Y0OjFQBs6gQAcDsjgIRIwwG0kQ/juSEsnNjQ3xYEAIoxBsGKeE/EnmZaKCABQzhXEH8MCUMMmACqxIkIwcJgPlMIpWudEgafmEBgcTi/x8sGEEUVJBHFUxBlz1QQSBQEAhf/MIXcoDGPxzJEEwK8SCm+AcqrlRBM+qnlK80UxoVsshjxIeQ67HkQVbZEJ5585oFcaQyE1KAf8ywIG+YhBf+0UqBxJOb8RRINQYyiUlgQhm6jIUb/MCBUCBTGwLZoZlmmcpmUoRjAgGnOUXlwwBsB6InUmhDuClBL44kAdFEyCH+QYlceFIZCFmlRv+R0o2oYQa13ME/8riEFpVAIGVoIAdEksczPnMDpkBmRPWTREYmgjDpzOY6DwlTgsSzHOa5Jz0FMgIZ8MEgHI3PTYNqEmuIM1xs+McGtLoeQ4p1I+YgCCX+oVAv5JM+K//9xwMMMgU+MKGmDvnoSGpqV1cC0iFkpYgUBcKiv/S0rOLS0QRD2hhUqvQf8WyrYzNakJSmdIkCWaJlD+KFSfQyFu08xDqTOpAVmqQEezWsBsOK2tWKixPzyewSKfuPZXghswqJ6wPYWo5aFpUgHhBVBU3J2oQkID9hxetwk0ufVbh2qfFZYj6hW9t/VGO61bWtQ8rBggsMxAWXmalyI6ja8JLXMQVggwIUAI1DYPSeUE1IPjf7DwBgtyD3PMZ7DeJUhyzRqV54rCdHW96F7NSVPhAJXgYcXgmA8R/i6EFcI0uQ/TJEAIR8K0Kqu579VuMQHBivglF7YK26SZMhJkz/Dp7QggJgYiTzpOckIIsQp+JXJFCN8ED6SxAVmPGZJ/4HE4Lajgz+lSFXJQhjH0JR9+EVuRNR7ETEGM/6FgSyFNZwVOdJW6dSeSEvnu0/nCrmMB8kn05dZTU+4Fo2kFY+1HygGF05jvAytEc3E0gdxRVNJ0OkqCnsgHzK0UocF2QZMRbIPKcMZi4fhJuGrsYkDM1NRlP6IIIWiDgFYAyBuPZGwv0xqA+yhjtPpM4mybOe/9LbgUAZNDmIxRQyPAkAlJO+kyiHFxitEBl/+bK5nq17qyxPTP+jln+pa6iTHR8OqvMfH0glnx/iZ8fgliAj+Acfrk1hplL3Hy0WCDej/8uQF6+ylV9ucTxbjAl+ghncwx42AD7AR4rcNMjKvje+G1htQpNZIGr4hyEAHmsv8LsxbEV0QwIgAIUr3IeSDEAkItEIifuCAL81YCnkU+R8czyiOI6rU6sN139MwRBUCEIsApHfy+x75AoxKaQx0dWCNAIQcYjZJeTQQBMQRk2FWmTHg+7KRpCc5LE2yMcF8oApzMASnfjHtRUdn6QTpOBKL0iEKVzOF+hcfQXUgEAcUNyRcEHoZmckoAdCozdsZASGsAQaRrDtB3RZJNsmyDLK8QC6I4TfJnWqSeP61rIfEOyOSeHZE79akxJkBgAvervtG9m9DyTCVofIEuO68v8Zk/nSAimnOTkwb8UXsH+kbwjnUHL07M414AXBdY5Hnnkwaz7M5aj7Q6wO8oFQmPHdJkggTj+RaE8wveYx9UJADxo1DYTZqTRlCwQCn3/4yNgPUcZc/xGMiTC+trO/rECUgfuQ91vpl19IwdkofNQqgPh/SaSJk++RhqwT0EdeSJgkRv2JpP0fqxbXpzVGyf1D8G0EZpVDNWDCA9xdQ1De3gHe64mEACCWYwTg2SHeARlfBAFaUYmW5eRfUFlgBJ7f65XcCExBOTBgQ+hdPgFACnrQ0ZFg1ZVDL0XY6hHEDa6fmbSaVj0bC23clQDhQHQdR41BD0DE0amBIeTgQfD/W+8xVUvFQgomhO/BVQrOgCEEwxTgmO+doAp6UMHxUwCAkg5uBKo4i1ZpSgSR2o2kk0DwXGPEzLVNxBS0FBNWXeWVn8gt3QjwQSzI3YS53ALy3gMEAhZ2ggFc2wIu3QL+W7bRIO8ZxD214C6kTxmaXf8h0MIhEM/BQ0PMToAJRKvgApwU2EOUQ0sBQRViXR6C3APwkhVOwfZ1Ah+owa1F4t/lgCLyofb9AxrwQlU9wAjMgBrEVTAYAhpYguOxYqzt16EBwC68TQX+hQMg0JzFhxCqkXyg2nwQHQJ1wT/A4V+IkkDogGSsXqzd4esBAQuogVOpYx4qw9LNgDGg4A5s/1/AUYG2hd8/AMEC7sAMjMAO0KDbDQQaoEEKUMIUzFW2yaIhGIIBZAAaKEQz6tMOoEAawEEa/AwtoIASZKM5URFBiORDKJMbBlWcrYd9gORw6QV4/YModUALdMCnScamCcQU6CK/6d4IuONBBN4/VKEaBENDzsD2/UMVoEEuONdAyOO/bd8uyKJBogEwSIIkVMEIuF22YSEaBAEw/AMwBANT4mC/sdUOFOBdbAjRmIkOPFEMuZ8i0ceITQkheSNhzFzHQcYSLEEJJIIftIAffJoftJoa1OEwIgTjxeBCvuNPDiIQlMMcat8xImUwAAMwGAJT+uNCBkPcSWXAHSQVWP/lLTRBFWwfFfjiP1ABQv4DGFxlZJKcGpwgTipdNfRSKwkA2wmEhlxiuBzAlGCSYXBj0OEFE7TAE+QCJSRnciZCLiTCIeRCLPBBVS2BCuRACcBj1W1hFlHY3qHgH0KdQEykeAaDJBTCFUiCMTggIxoiQQQcMlYBMCADMghEa36lQKhmFRiAJAyEfSrdCLSCJQSfI0xYbFLXUpHDLpBhBHGAa+UUkynAWT1EAdxfeSkfx9FITbUCJdTitZniHf7btSVZQUwBUBqRZr5iLFRBIPxnPvpiFQxBIRRCE/zDLVih0tXhQaBBFVDBEDTBLdyCDZABGAwBQVDBi1bBQOxnQMb/mtvxgiUookCIWR7tQGSOgYJCUE75GOEV0EmKFWOwJG9mkkAsQSLwAqw1xBQcJpIdBBBMQZsORAxCZhU8Q40a5GlKgo/23RZem+shpY7yqI/2wUD0wS1Ign0iJBnMaJ0aajAIpNulgAFQQS0uHRD05EIawjIS4JU+0CwwkAbSn9kBHUSIo2FxAS/kwr8hxNGJwxBEZg6k6kG85j/sAK0GQ402QQrs6Ffi6T8Iap0KRB9UwRby4UQiqWqGZo/+6oaMQR9YJVIawBDsJ0HcgjgAw0QGw2mmgMnFnSPg6AwwnSFcWxWMgahKkIOGqUlYACFZVGNsHPL9GC9QQk/+G6zG/9SbPMMOuGOAwVSDDYTrjWaMFgIdFARYDIdB3II7bMgzBAIKuh1+okFoksGP9kEfdEMfjMECYMMY1KkikIG0CkQT9AFMUGvABUEGfOW2XltsdkIrzAAfUMEMgQOYoitEIBQDsd12uGWMCF8LcAEXtEBVFcQcTcYcsqhAeFC/FpvwPAQZLAAP2MECMKzb6SgaWKUkTGwfuEMTGKxAQEE8xENCgEUMwCdYDgEJZMB9ZuEOzFUQGEIrBEMwDJOPNEC50uxI3AwmmCICDdV81K0C8WAC/Vua/kPCEkRLBUEtKgQ53AJYUAQc2ME3xEAgBIMxwGe0hmzWXuwCxIC/GMQqKP9EOIwBfO4nGJxnav5DJ4jlHEKkFpbDDuzCMBFTYP2DcNotLNmuWH3azwpEtlHCt6apJRTECc7A0/XpQAyoCh7lP4ACQtCtHdgBLjzvCVDAuP4Cs4aAO4yC09qBJVKEEogDfbZmtHalasoiFZxcCgBcK7SCQDyDQHgOBVJEp81Hp+Lu+nmgmazTlv6DcPEC+6bpDMzQERSEMYxAJ7QTWRrdCJDD4hSEjBbEoECOBNsBHBQND2hvDHAvfsTOecCBhtToFTSBJHjsfTYqwGXraf5DEDgYCniOQMSv/cawfljolLBCFBjE6HHBPsjrCHCmJVCBZRqEJEzm4yHEDqRc6yT/xNtQDH64sNrhx8ugTvc2xM/oQgR4SB80wRAYgLH6YhBQQfr+QwqkwNONwBikwTf8A6kIhJUIhBWYx5AZxuhdYjVynCQdRPzpx5hklUCQI/+SES8AwxDwQgakwD5kQAbwQhgPBGlepUEC3Lf620JWrmQsEBnYwi3YAhkYwECsMBCfrEAsYTnkgDHEwRrQbSAKxIBORJslxAEYXmHMMSOlwR23SMZ1nMQxWy1AhhPPxxEihClNAAMQgWz+A/ECwwqv8EKcr2oqrxrsgDHcAjmYBAGBRjXT6NZysgp/cUQucicU5j8Ywy+ccqhMBBuYAie0siv7ph1/3pR4YkKUwRLw//GJLUtfuc8sJMIv/0MrnNxBiI1BnG8GDEEKiEOA4mQgIKlhXLNj3MIfQGoKU4EByAMwnGYKnyA0B4IuoDJhfBVEsDMsi4Qs6yA4/kNJIwQ9C0RuDsTMhotwEQJCsGED1S9B8AIxhqcyR+pCcPKdguwfoKdAGoP7/sJuMvRGPC8P6MLT/gUZkEAhfOUXp0AG6HTjLWQPGIMqoLKM0EISJe1DLML+KgQ7i0IoyDBE1LFJG5YIGoRMS9As2DSIUkHweqUyKwQyRCuvKuotUEAuBEIgkAOc2MHLEAYo9XJCTHHpksEWp2ZEEmmOjoAjqIExuMMpNxEtKINXO8QzhbVZN/8GWoeXGr5R2cE11KXwQ1hmBmTBEIxBDOxmviwAOWDFGHwD5Az2QLgORDzv+zqE/AixJEx1RKJtRR9EFi6kChDCOKMyhgAnRJjCuXY2aNxyu1IEFzFSSztGKb11CRRoXQuENhOEMvenGH+Ch9w2OPBADIzCL+iCUZvJ+aYvIjeEITCsGqTcRoNgQawyQ3i0DJdASivQdUcUHHzJiTAAA3ABBwDjG6vwTne3dyuEu8RLe+tH99LK+X6lAXhlCgeBgzO49skmC4xBZYcMdI/Ef5e4QvBtQpwWfeQUGc1CCiRu04H3QSQzVDt44aZP+rAC5EwxhVOfEBSCY9e1aXc4g5//XCf8rhogN93GBYpDhBqUEIsn0OxehukNRB5fyRKp+AHNAgPMwiHo4j8Eb0IY+X2K1fmeINMZAw80wC/kkRUsgRUsOAO51vQlRC5Uwj9w1wShms260hrAMEJA0rtOybfxY5dzwFvrYqYihHgPF5LPQLcucBzQggrwMZ0HXUhDkXTrh4zcAc066Cz4QVaOuUE8+oB1gpqnnC9EgTyXwZxn9pOLtkJUN7rOAhf84QicZhAEA5kzeIYvhIYTBKqbSbFTxHCPuarXYSwU8E1llRXUqwQ9AlrOOkGsdSqJaAHherYV5AwFAS94+ENYNDJ/tysFwQmqQXIi2w+ZSiUXxJSb//Vzo7iXz8Is5EJACgT7dkK4hzsnf3dd27gnd7KZg4bQKLR4e7K5m8TJBcG3qkEnWEIZlEGmHjoL5cIc8bm1T8Qc3fCNfAAHQ4S2F8RLGgYIxLuA/cMsJDgLqEBVtcIIUEK4E/s/LDxUn27N13wQBHsKz2dh4AcPQM7UMPjOn/l89PoJUkIl8MESLOMx0PDG50eni8o+KwT+FgbP+O1BYFRQOsSJi4T6MQQXIAAw1ncuVJUh+LsBHLt3AzEwVKs4VMFVikM43IA4FMfPf4VA3P0NWAcZBDHbgwYaLOQM+O4IWEEOYALUR/16kOQ/yEI2WcO7y8dNNlPVm0k2etDII/8EE3D9RsBB2Nf6ZhBCLgyjFTgegIKlQCwyfwqEZRKAEFQAJPyAAA3EgiTPSNAJO/SDE2ANPegB8OuBMLgC19JHXYcrTO0BJSxB4gtEgDM+sVHENhBEoZMeePm4efBRLlgCC8zA6WObJRjAvxfEo2OBFETDO7wDaHTuQIQDPUTPQGyBX4j7enzlo89AIFDpHjzBWALEP4EDCRY0eBBhQoULGTZ0+BBiRIkTKU6MJZBJRY0bOS4U1ZHDQE/iYo0YMePfjE4pgDWkgORfs44bV8zUaGnElH98Yr2Js8ZmUKFDiRY12vGJQaAKkx51mnAc0Rducs2wYvKfIQMGEHIVKI7/QhIp9J4urEEwyL+0Zf/xEhgkiKFAU3awMPZrzT22e4ti0cSXbw+DGR9yYNBQRkE8BH0BntnAcUI2AgNFOZRridV/rVIYSCHQq8EhZGrqiXzaIZWc/0Z4ohEnDBGEUlAfjFIbd26CExYWK4hIt8I7FCEv/XcNtSmBZ17kopR5iUlLXMUNDM0V2OgVZIN3F0hlhs5/ns54X3ihqdF2/zQY9EFUvMZJ/47t5f1PuXKFkAteEPhGIAB2qO2ixCYCCihATgtJoNvu4IWPGZYQKBdePiNoCEm8kuSfQpwwT7e0qPgumBHK+YcFt3jpwI+BTvhnGtyM+4cwgSoB0aEABAIi/7caBUrPocMW4uOgHQD4BxPcDKRoRgGWiYyTRf4pzwJLKJmBBdaCsaSzgYYwaIUxBOLhnxj4golMgdwhqqV/rjvowoQMiZCucmagpC2BIBkIhH+4CK7GEnB8aMBBGWKDQUNP8+KBJyMDwYJYEuHjpH9iWelLRtj5w6AI9swtzaBCEyoYNGYY4Z8dRkjkEB3WgAMdCwTrbg+K4kBB0Vz/mWWgRHUF7IGBuInMgg8sYUGzNnNNQphTdB1xoFJLNUnVGYIxZgQ1BprnH24j28PHiapTKKpfzTUqgVeeuvFcgWQVB9t/PhzITEU1qfegH5x9aFSb+v0HjYAFRimQWHLhYv8VUbj1VqD2GETnqBtr/SeXhuIYtqJyEQKw3Zkm6xgiHv/hLZGOLQCBECJCQegXjmACLJVPUzEUDSpqpiIINEoMJpdtVknnHx800OCVP42BmC12GzpyKACrARlqjgqNmiIKWv5nAaoJisA7NBAakQqcp+PFACoMGSGWQxC4gg5QeP0nGxw5fuiAf+puCFWt9T5Kto5fIOjqvcf8h4eZDYXWzSC2MgCYFMRJoZNWZpiBD15aOORqvYbyb+KC2nkvKI0VSlLwgVQgyILSy5rPqDL+WRIifBPiWvWuKIozzoW8Vgu0znxPoTMDDDl1BD4IICdwoSouyIf31pvp7oaKGBT/AYEGoEiF1GtX6ILO5dtecK7+hSh3iVryDHj0fbeklZNGMOQDIeAQSHOiQAd/o+uFhOh0hnzFLQHeYR2InPEU2QVnfP/40l6UBTwHOtAzvAAPtmaQCwwYzikauB/+InKfimhvIC0QyCJMsQhOPGQP/qFRfDYCDxN0wQQz8Z7F0lAQLxiKazl0RgQKaBQexIBMoXKKEcyVgiEY8YEOtMTk0MaLZ6wBQRKJgtLKUjfRgUx/AvFgR1wQkRnOJIa1iUMNddXDgejwH2YUCg/8MZA2PuRlE0lgRBZIFCP+IwNIzOMegSdBJlKiCtnQAQEaAhnI4IKDHZkeQqQkkP0JpZEM/6nVxLTVEROEsSJAGlQrZkK7M6oxKGnSF+EGgsGFZO2N/8BGQyBgqDh9iY8ZGEIsjci+k7RCHIEgyAm7eMJP/WNGd6jEFzPInkRy5H+A6UICukARZRBkeRJpxD/iwBYZSKAjntxLHxZiBDCw4x9gUERBiDjOicBSIZ+p414y0M5ZtjMFfDRAMCbHhyEwgxkC6eI/pEQASKwhDdW8Bi0UYoL25OqZTCMI6QaSt2Maiore8Y9/YMeRrGUNlEIBQ0JIcZBPkMIIRNxL+TIQkTjN0SCfaSc8VxpPI/ICDcVrxT5OyIHJuMCm/myAKnbRJyQNpAD/mNgsZFHMj3CEdQp96P+5bhRNiRoEmxzh2gG7A1KRPiUFWSjfP7LAl5V+NY9HTIHk7pRPTmyADS4wBRsIkIoGAKUxO9iBCp6QCEq0wHIt0MYw2lO36AVlgzY50iI5QliKiEwj2pubUzC51NJ9IpxEhCxBSNHRgXy0spk1Skk1stWtKgSWWXinaMHKi05UCp9s4ASi2EAEFNTiFyggByEOcQhetIKsTGgBJaABtS8gBLEQMWxtLJCk4ToWuR2xwzecYU6B2IIH2HBGNxQBBsiKM6RG+MQfnLEOm3Q1OF3NQgZEO97xyrKdBuADkXjBC0vYtr2UsFInmHiqyU3urnhCxTAaZi48/Pa3QQlubRb/m1wDUwSRAnmELcYZUu7+wx/veMcj/OGMmnyiurZwxiNUyRHwCoSzQVnnQUYsEPOSF8XnbaclvGYI91IuJTMowX1pLKE7teBGJWOLumwSYIH0L7ECOW5BrseQY2DCxxBhKIh0/J8lH9ghMcjoRhL8j3WMk1P/6MY/ODzhCWPjEdJdwCrf8dAsnBnNKUbxEoOBp1YQiZ73PckMYrHemVLiAirkixxYWJEv7IIgOYByZA7BFkcFRc8XCJdR6uUMqlKEw/54RAyy/A9F2ALMAynzhB/xCERm+ikhlkhJS9yQrpL3zKg+MXg7QU+3pCRCweCDISjR3gzwggu8wBNfhDaQ/yFTBMC/PsoNBq23RJfF0fSaySoV7F0sj+EbHEZkpCHMYQqX+Skf5gt4j5AFeaAZzSaWBy/m5DV+ZGAfK5WHO/mxjVwQSSB6ZktjKeJTPpUlkg0ZoEGSLCXl5PtcbxCQUQ59kJUpQFdcmzKkB/KIb3BZILjoNMQjHWaCcPghtziIqM1zhH8cAeRZ6Ha3z4xHPKZgTnzYx8ozsI2VntsY1QiEDOQtOBAKRFAD2bdRBCCREgL8IZoEzNOOEqyFrEw3C6CNoiwuFG0nxOMe54s8jkB1kFu924X4x7fH3YlZp+Dc2zgCP3hhDIFMLSgc4MRagzMh1hxWI0rlN0Hy/ciG6P8Z7aVThqMaZXDH5FxrGJ9IEyayDYGI4SDIKAjiP76RqH8c5CMP+be7Dbk5pYAZlohPgYsNkWk+xYRBP7AjGIJ0jsjhH3Io9ECSLBB4CwRoBVn6QBZelirbxAYEebpApI6QNhiE8QRRvOI1gngxHOH4yY981UG+DQnyAQ2d4EIuAjG1N6gABv8Q+kSq55CPILzzNqk5YG7ec6IA+SD7LAgXbtORviVk+zhiNl8er5vjf1z5xwe5/rexj1zImg9aAa9i4WnewAJYIKiCSiD4iyAOSiCeLPz2Jv6Crk96TgAEgOh0ozw2woNaryAUMAILovcaryL4wSaMDxnEoA3E4Pj/2iDyjo8f9kF40KAV0IAPao0X3o0PcuECcuEJOuAfhuEj+EsUhqGoUqUA864hRMcBQ5Agksko7I4ilJAoosoJo2YEJeL3iG8jVPAffu8fxAAZkO8I2iALYBD5SsoQcGtO3qxkWgAOeYFX4uEV4iEeZOEV8nAVcoEP/cDsOEL9QnCLuu8KB0LQnqk2Wu/10qEO/yEqskYgILEQCwIMy2ILBaIN+KENkGEFV3AMWVD/8mjX1vACWqEp1msHnUMV3y0WWjEXYoEKJ1Ej/kQWdQPJzO8fzE8GDCRdHOAVxkEEBkIHsGZ2/kGboKyVgkLrEm8gFK8S/2H4xJAFl08exs0S/3IhcrwGt7aRG7cxFtzAEnQpA2txFgmCEMgxKBZtIXYBAPDgAgVABVhABkqgruagC/DQAeYhGB+Ch66QCyVCHngvCzGxlSDgGSHAGTGRH8YwBf8RxAQiB83GEAyBCjqBCuSLF5gBFv8jF0OwyNAR9AoiEBcC8CLCHS/QAkagBOjxEOzRAbqADqFgILKmAo4x/BxyJj4sIA2iDQyyILjQBCkRGnlP+SKP6o7yCMSOH0DBBMRB7iriCPVmAD6SAkDSMRZhJGfiDf4rFwXAAnKgBOSxABTAAV7yJeNhHnBgIOLICR0yGUmgKJzRIFsJFOASJ4fSGTtRDJFvGvmBL4+gEP8gYBXo0CoL0ymwIP0cQgVKQAYm0CDeQABO8h8sQALCEgY+IBSY6RV88RXoIB7Wshbdsm3gkih+DwIQEgJIYDSvwCAM8vdeUxpT0C/9EhmuIA/ygDB57BwNsyB0hDchwgoPwgMcIjgf0CFwZSCwSQJYADPnwATmgA5Wwd2GYBUIrzBZ8x/ogA5IcygSciBaaTS5EBlOEzU5cRqPTzBBYQ7ioSx57B/cEx2JAPUOwjcj4R/I6DcTAlU8cCKiqgdeQNgGAlfwYDH+AUBYQCULYB+2gRlyLQBb4WCwcxIr8S2RgQRAYTuTMSjEEy9TUzv/4TSvACGRgR8ggB9WAUVXIQb/hyAXzjEB8uA9C+KE8vMffFMg7PPAZiX7OOIidjQoTmdWrOcfPpL17K3naNFyKGHXNqMVDKHOggEZDG9C/4E131IgbLNtBII7nYIErgBD50E7SSBKWdQYBqSnesANLiI4nlJX3o8gbPTAviBIJwIABO4fAO0f7iBLgmLIZEMOBkAcBuBPCSAKUAAFLoEdIXMHciEFgopIHrQb0YBDcIAtJTEyHo0geshSn4ILVRMUCmIVCmJLh3IiWgkuSSA1ryBKtYEXYPENXvUNQCAKLiIX3BQ18BRPaXQjEiErI6NA/+FX90JQB8APANUPCMATUAAE8AAFTlJVekBNVy4FIJUz/7LA8OigYyqAGBdiE0pVIDR0IE41O/PhU7UQL891IcQVLm+NC/ahQcVhBAJBBYwhSzjhOXFDoY5ETXNlNwFjTzliR6V0Jv5GI3bhV4M0ClSATSuCsFrED/5UDuQAWUEABHZhFy4QAALBGPhwCHJtG+WrpNZt6xJi9mySI/DF0dTIZGdyWzXiLslzSzWUNEEBQ8v1IEbVIIavIbiwSv+BH8SAF4ChYnhhH2ahQbnA8AKIIPaRLQy2EAWgMcKvMYaDL1okYiU2CqKACzoW1+KLEiaSDzrBEtopIA2vEHayINiydloJGe7yZlMTXA2CZvMhS212IEI1ZxdCQm82XE9z3f/cKxeusb1mgRe2QRsUAPwGwgI7sihw8QrhVFcC4BJMhyjaryzkk1DxwBjaKxcSoUJ4gWypzttGtqvQdhmXcXsKgQ4KwVMFwm3BtSBRdSEw9ENtgjVH9QpOVUTJ00TPLQMs4RqtxBKIwGfm4E0Z1ztogChs1TBx1CnuYE6fQvUK9Q0CQRzkawj8ciA57h9ugALCQRzIgGlBxAwUotIEoipzjyDIsy5Z023D9R9OlQTmd34PAkazEwrooBfstiK4U1zhFlVRdRV4lx/4oTOosyCGsyMd1ztQQHmDtSw+oDYs1zwgsCKQ8yHmkyGOhD8Nog4M1WKtd5YIIiBxwAYw4C//YqKAzuEfKoA2kqA7YOEfzmIgzMAJCkHbpI74VHVEXdeHQYEMtmE7/xFve/Zm6bcuSXNUaZdu7/dK15dtCQJntVRL5xeARfQKpFOWOCEUFGAVFGBvC2JyI1At/4GQ/oEClMAxNlBXI0KCCYIGaOASLiEACOFLFhIwXUEY0ightLU7aFggBmEQ+sHwPqz+nBHxytALSRUZQGEIAmEIaDaMG4J+L9SS6/IfQOF+SSAPaDd/28Zmt7QSJVSJKxmA4VY622365IAT8PYfTK8jYHlviBQhGsGWj0KXfsWn8AByjeKMh+ISGsMXJjd1PKEKxMEDPMAV/BiUWHiGCUJMBCKa/58CkA1ikMWOBNH28FgwDDexDS6R+EBhG8hBAJ5BiFG0NeW2IOqSnWn2Qt35U+NZIOggD7QBRdUTFFC0lXa3S0lgFQJ4fnP3nd2ZDKrgVWWlB5g3lvUGA5zCGgYCghciao2CGiZCQYCVTzBYR8bYPJw3RyCaIKhhBfx4IJx5L6qZIGRYIahhH0dQZxcPGjdxLl9znsVhF3zhDcwZOr8VIfg3XNn5koP6NuegCpgjEFDgqHcBBZ6BEKpSHMQBB3xmFZ4TjEOBE7aBEMjBUGvUcaM3BPsVA7CgXw+ioSvioWsUInyh5wi2/ZQ3N7xBINyxdqK2FhKC2HCgJmRiIJqhBv9qYiD6wSZQ+h/0QA+aQa//QaUTwhU8ADu1biEHAvFckAQHoifHczzJ8x9WARTCIYRR4AwIAQdWITrzObMpGajzYBVuMx7yIAGk9G9eoE9QIAA82jcDoQr+4bYJ6Zchd6IhIqIfCjEXoqw5wjcn1xsU5Kz/oa5rdLlxZJoCQEd6+ZiqEgdcAQcyoQJ+QCAqgB78uigI+xxkQibU6Ae0VbAHghr6IRS2YRueWhykGhqPIAUJAgx70r5Ps0vJEzqHQKuZ4wyQWmPFIRRAIR608zb5t2b/ATc98zavYF4Eog6A1d4GwqPb2CbGeiKcF0cnt5r+4aIHohiamyDU2CCSxyn/FAQQKrxjysMTKGI+q3uPDVsYaqAG6IEe9GAQ/iHHKaLG18GwtZuPKyLHqQED1FgAhAALMIAQtmEO7BIaF1JnexJEKxu/+Vm0cRsFlEAJxsAXfGEXouAZlPyph2AItoEMhuCp/4EQnuEZKKB6qqeiFZgiwmCsMbwgelshfMPC2YLEDwI4CCK4jeLDg0KNY/tXbsB7W7iFZYI2mqGiB2EFBFnHB0KGd1wgZLgGhIGkzeiwM+qwCaIZnKEZkqAGYGEQXGEQAFkJwgALkhwLQpsRRJQnQRRE8fuU/RlVWXucZdsXauEMWl2sCUGCMcA1/mFyOfofyhgh/mbCGSIMyBEF/xrjt/HnzwUi0IsCEOJg0IViGDWiwydCCCDCFQTCFVKYhc9BGMLBFUY6JlqYHroBFmTY1BG7G+ihArTVjEDp0yFCryugBlxhC7y721k9DDCgCpSdShGS1mu9IG89d1P1QvOADJ5hciNczZ/92ROCDASC2GwCCzIeuao9OL59I/DzeN26ISx+KPR8ILa9IEyeInKZKJBjIVRBIET8IFyBAnAAA0xjj10hE9rdIA67AkwjUwVi34dijwlCEAaC1TGEE2zzRTX7n7PY6vFbswdak6VTHEic4IMb5I29I1RcIZA9kWCrO+bnKXQA5RMJgzuC5AkiDnD+IGiB5RfCFdZ93P/3PelL2jH2uAZMmu4FIhwO4qkp4AzIoc2rgACOuQowIMyfAQueoTxyGboVQuY3YnLJ3jHC/R/WBMJRw+YPYhi7fc9tAua9Iw5o/h8ISiOqEugNYoX/waRrHyFIWiBm/+gVAvcLYukVYri7dyCIbQsCJwBqIQCKIQB8IcQFFFe2OiHKo881/x+SOzciPOx1Ve2PKfVRI+4FoobSADlowfoVAuXrAANWgAJEWtMPooDMyKRBnfYLwhlIuvdzXyPu3yUMohgAolixf7UE1qr1T0fChf8INnwI8aHAiBQrVmxkMaPGjRuFnKmIgqPIkSRLmjz5sEGDNQ/hPEyDsqGqmDT/a1JUYjPnyVqXFD4M92+FsHURz+k0CtEZxArNUNL7l0RkHZEIGyK8WouGxao6u3qtSOtrTF//ZkI0KzZtw5VrXP5j6bYBR64y/6VKpdYiWppSHircGzNT3ohcT2z5l4kevagNidpUSrFp5IeSOVb4N0iPnn+OtcZE2GgiRoiItJ7453mwydSDw6omaU3mNbt5Nf0T5FUlRJYnEUF6qMqsrn/DX3vt2xfiaJO41XL7B470iVFmVmh0XPMyRe016a2w/pCeKyEmt7j7lw2j+oexGyKiSMu18dkRfxl/iPH9/f0iydtGoppcg52gkE/8mQTIP8tx1BxiJbkl0nMUNfFP/w0NMQaRMP9wd6Bl2mH4DxIrYHDCaf+Q15BgDv5z2Ekn6NchIAkm+A8g7VFkIn0ZYfDQFipG1AgtowEW0W+H/RgTjBbR+A86g/1W4Gu8vSaFgRnZ1mFD2TSUIJEj6dgVN3E8hA467uDQzUYVaJgTh5xZhJRIRIEHUZoU/JNcRYIhmREtsXnJn5I00mfiP6cVChGYDbXYUIMUAeKnRj41+NRJNyKHZ0RMZslpToiW9dBvEKFoHA8RXaMKIIBWhCVNEHJkB3ThiGCGDUlEleZDmzyEnVduNvSrmkmsYFsF6xwrzLDVsUnRrg0BqFGC7YlakpI50bdpQ4W+CJGTNVKkSf+rGm2JnnxfKUpLnhVlu5G5JZ2ibqcaFZcXtF9F09ApkEQgqqizKapRcuTZm5Yd4TBiw0MhXJiRMMFmqR2zvUL1jzAruJIJxv9EkOFDwpDKkSr2kQQjuyKlMtMveKnlbE4RcJxTNoCgsypJMP9DbUZWyksTKw3BxFe8IwH9z6sZ4UtbBHehZK/QNr06yj+KmLQOs/I6xqzVESWLsWAUvEyTk2jVDByoMeXM833YZnQzSdSmYjJ5OoBcUWVpVxTNmHBIE9PKTmcUB154+VwS3w+tDBHiGzVlt1gxODE1RAnTWVESaWI48X4VDFvDmhuFAEYyQCVBwQpKL1ATOIpz9Bv/2RqxIjjhd3e1upPXAIxzRRJq9JupqYxp0d8Q8SA4D6c0xEo0RHeK73O4eBXBDw358/zxDdH7c1f0RrdR22Kt1ADoD/3REPlmjMRIMop0s0DLbwI7mB4XWwdiQ7s6lg8pyZjRzWIZIyG9hyilcRXh3piwB5EYPMQf/whgV2RnEuDZhHvEMdXG8iWSpqDtH8/xGeJYwQ1IQOIHp3AgRHQBNMNZBIIQQY4zhNcQXDziH9LwmfVmx5LiGK0mxzve835YtIakIg0+e572KIIvFZ5khxr5xj94YIPzRYR8QMlVRtgBkXwwAnLhWBifKCaWJITDDIOoWEM0tKskhMAJUOhFykPy4YQVZKIG9KiBK2ogquiVRBcIPOE/TuGPVJhqgx2SnQRjQkHEmVAjMINMRQhHxH/4rHcWiUNxkGaTRWbEiLOjyDROEg1ORgRxuCglJFFIQxbaBCZjSgMQh4MLVaalAVEj38L+YYt/JAwoELFQRKKyRkZkMSKMIAUjwLAC91WkG1YcSRIs5ArKEUWMWHzjP/LxD2q4oiH0yEQSomm3G4okVhSRZSf/kcK6iUQXhxze6hrYkB/wqyFNOYU0cGE0S2bPcAzMiTkTGBAAIfkEBQoA/wAsAAAAAOsBGQFACP8A/wkcSLCgwYMIEypcOPDevwYD66UZeIygtzgCAzDcyLGjx4KLPoocSVLhmpIoO0JkyCJHypcJJ8CcSbOmzZs4S6r4JyGnz59Ag9Z0KLSo0aNIUU5MyrSpU4YdOvyTKlVgIF8olAwM9M+Csh3VBAIwWA7Tm387uEYhNIALNAUJBCp4SlfkBA5c6uodiYCksoHS9tKVAUOwTXX/FHBJxGLKwGpeCk4qJzCyZaFTSjyJ5dKnjH9lCp4VqMswU6JOL1RS2KUp6oMCPJ40TdtmjicuFMyB5keFl8gH/5I9Vs7L2NgeKQtUjjLypGpTcuXFyeLfGzyjay+UcUF73VDeBa7/DF8T/D/EMIksxPSPD59/lCkLT6isohdlwAsS94LpGPt/YRm0zEH5DaTMgJUtVNEkB2FyCANMTUfehE3Ntdc3A81G4YbZCGRMQcwNFOIDI/CRiyVVqPGPF+UgiNMD8P3VYov/YIJJZOyxVw0m8Q0EwFhvjBVAAJEEgAcBnPzEAIRISdjRBd3tUZCGG5JUgHasGAQIlQNFURNyCDk0WyRj0aSFBGX+5AdCxqiwA0OOwVeOMicGE+dy8NH013wgCqQMcyHOx6eIBgEQiCrjVakQkyEp6qhH9TwqaUmqLGCMYyr+A4SB9E1B4gx5FiToP4OOKlAsUyjzwKD/PMDcnVOM/2AIGh+2mieMsRIEI0O7/MLlpAM1ilM7wBZrLFNroNDTP0wg1EIHHxijRmdqjHCnQZv62Wqqth40Qi6xUEZiMIb8E8gM5QpkgCRVjADiuQKNUM4bgQQzkCQC3fIPMFUYYswOwaCRQhaFSGLnFNkWtCtBLEQRyC4P7wLxPwv8A4c3x9YVV8Ycd5zQGNX9I8OVLeSy00Cd/bPTySygquIUMB+kghrcbuoYjB/2EcItwQRSLr6KNEFQCAL1UYUxgcAoa7oCATPEP/oSNEY3fUiyLhX4/tPHQH8AM0Igjs1gSQr/zGDtQGpwlW4wbJOTBpcnV5lkkh4VdgZMsxRkwj97e//s998GMTlQLtXyYYm7xmxDDg8xYFBFILJS8Y+9/9y5UxXP3IIBGMkglEdB9uBixz88kC56DE3cMsYYWxO9tUALhPPPOBthY8Y/owj9TyFDICOJJFQEMYK7lhhiyb49OzYF2IEE0sQCv1JoiuA1EQv49YbdIVjeDGzDCyWddGIIMAYMkUIKBhgwkC2670sQMFRQEYy7aqgYy0Gl1ZW/QJIMYYDk//ifATIwBPL943gqW0ADIDKNgXyjFgfRwhewlzFKHKUEBLkEBSc1AVP8gwGz4MXw1BCMIBgAGANBIUGCkBAIXGEIfViA62LAg1+MwR02CMcCRgcTHv4jSyUZQhb/1JeFDJiQhQUJAhXKZYwTLNAeD9mgFPUCxZcsa4obgUdKZnE4s7XCEgawRPwCmBAkFkSFC8GFQEr3KGCgYQQ9GAMc7rHARI2EDSTxAUnY4IJ/sIEDfbleYEqSpgk9oQSF2VARNPWPRdKGE7NgjNliQQlKjGAGnUDfP3ixRPWRUV1YHIj64De8WChhDXVUxR1KgMF/LCGUTYkAQ7gxEDzAEiYOKMU/dJmTZTnSMFgghDj4MINiXrJsfEjf0wyyzBSK4x9bGIUUFlABPeiBHnoQxjWvKbuXbEIgjHACDm5gBhuYgQw4EIcBzFgTFAJDeCNQgyl1kQoUoAAEIFBB3G75/xJi0AQckSiJLfmpnQkmZQPDnEEZiikQFhiCF+YbSAqaKRCyiQMJzdgmPYCyUYF0lCAUwIFB0HgTQ8QzniX43gX2AKUSSEAA6FgDK5aypkm9h6AikZKUOJIkDwoEjx7pDk5pQj02sGEffGjFDJSKwRkEYR8TXUjFhipK+VlhBlYYAQtaUAkW7CINDUBlBNjSgQmY1Q8TGAABIAERGghEDlSNq1xRYj2RooQDbGCAH9wzg1iMgAvbYIgsJaXGhJwPJkGYn9mGN4JYEIAIE2iBWSeAVj9gQRoLpMUuosCFYWjgAKAN7QH0yIDVKAoaJXnTm4Lyy5r04B8v8JIF5nqTA//8w7YjqalA5sYFN1DiELHIxRVgh5TB1oZsBEHuR55mgE7Mz1pTcATMplAOmNWvZbngxSpWkY50aEAUPhDFKxbjBicuEJWotGOVcCuYhBVlAxxpxVN8KpCz/Ge2HZPJqYap3awRRAoUu4ks2ViQBRiYIaPY2uuC0swMdMTBBWGuQVioQrJZOIyzKuZSNRwLYxoiF6PQxQngOhAX0O0gcPgHCgZi2kkNFCUvSAp9PSJftKSFtjWxgAVUwItc8OGZ/xhDU7rZDdYpghRGMMInbOGMJndDEQIxQkE+8QcnGKUQH4GwYTeShSwQxMH74IUhlvoPpVJiG9pgxh/FAYI3+ML/F3iwwA70yYIlVIcPZXiCNkgCX4GgAscH6eM/OHBiQNPlC/i0wBcCQYkWvGcVRINJYTmCjX/44xHveMQPwsEOMKxxIJf+xyP+8Y5/TFo78hAIln+CZXlkYR/FmwEaWtEKSoRZqUolZitKkNR9tKAFCBmGd/ALaFOwQVgIcYBAtKiQXBjFEd1CiIVychYQFOQJ/2i0JbiwiiCHp9IeicFL+PGPIwxEDBxpw0FSTRNzD+QIR5BHvI+QBXpvQx7yQB8VOkFr9/DBEJ2whCX2AVjAruIV5IlxlYRFPYR8RjVCDWUhi7ILhwukBdDYhyEKcQV3IEEI/wB5QWRpXJyq+yfs/x4IMv6h7parfOUwF8gRxDDzmtMc3kcoRLxXAYp0xGMcoviuBkohCk70ABM7eIPSbxnIhIBpfzRplk10KQpDK4QXnOQFMwi2jUKQIA+Z+CYSrL4QCOTk5N0GxSq4MAQEIIATDOAEFxDABULQS+l4f4MFYnGBXBQgEdCQRSm+KwoHjMMBrelIw/kJ9ZnIwA11Ceg/wESbRrxEYvSygDGeQIknVGGT//5HBuRd7ywg43MziYFxndER1nukAkchQT5AIRAS2F4gZhfJyj1idgiQAALAXwXw5RFmYFhCHLwg+D6WzwVmhCIPc3hFXFBP9urTxqD1rTgB/sEJaISCGdrYxv82hiCOE1HCEsknPb0LQbD2w3t3AykEFDoy1aAA2Ca7TwkJ/pEHOsw/D/v3D7RHEAHoE/u3Cm2ADClwPLzABbMwAKFgIV2QABtDHta2QV7SA1HwWlxRcQxBYhe4IXfwWi9wNy8BAAJQcRrxD9v3D3JABCSmBG4lTEMwBIUQWFewCsiwClfgCrDHes1wDgTBerAnEN/0EzWQELBAEEtYEOzmbgiBbgLRcnkwBGQQfcDne76HezeRB3mQDwMBBXRAB6AACrYHAd3WbWYnfP+wf6DwCmMYCk4wBHLwAWeAB7vgC7uAhymIBy9gAYHwAeZhEDdwEC/mKHhwiHURB4DwD8X/QBAQxBC14FYp0XQLIXn/oAoFoUH/8GK0IBgasYIv4SXU8A81EISupwdJMAiDYBDUwA4pkYQCkQRJAHvN0AwJsQL/oIuuuAJjEAxXAAFHsA3IMHMsp25SqBAQ0AYQAArbIDEoEAjRKBDPQABDcAXQkAdv+A9keBADSAfcmAdwOH//kAB54AEDoXAGEVCY+A9YgAEGgQU6EAAeaH3aQYkI8QuIIBTsKHmNOBAYsxdLYRCWVxMh5QrCUAEVIIT/sIoroJBFKBALuZDrYIpLWAP0IIS4mBCutxFNxpD/wJDnkISZ8A+CIBArJhDvyIL/cAM34AFX4IX8B4C0l3sEkXu///cPB7cKOHAVEKQEWOCO/wCPA+EL/xCJAkGUBXE7BGGC2FMLjxgUnGgUKwEHg2QTJYcU6PAP19CIgAAIGOERxfCJjggUA1kQJ3ACAwFgW5kQWkEBK0BOvPgRFZkQIFkTsLcCSSgMdTkQmiAStPCIZCkQEISPAmGYBVEHdPGXDKGUAkEBBgFBSGkagykQv8ARankCEaCWNRE9COGZ4XENmggOYfkRlzkQqoAOp7kQW3CSAiFyNQFEYfmJv5AJZrACJSmLAiEMM8GbPlEB2mQQFIAIAIYE0yQQjDkQW/APH2UQHZKJbTkQiPALn/icH7GcQykQ2PkSAKYDmfgRukkSnP+ZCbq4nOFZEOhgDXoBCZBgjxviQyMhZEtpBuHQDQiRBA1Ji/9whE+xDrzJlwSBn//Am0lQA92ki8k5EBHpHZCQCv/goA56PaX5D+BwEJz5D/v4D6UBRD/RQFPyD6D5GiMxHuo1EhiCED8wEKfAoRp6lhqqCyn2oQzxCNFwagWBC9EwakLRACsAZQahCN3EEEnQo8nQC//QOb2QD71ACuxACv/QC+wQDuuQBH15EFQqoBvBmzWgi4OApf/QDf3QOckABWCYDMlgAyuwAmbgCjVQoPbZUSnaEYOkRqwgDbhwlanQnv9wCgUxOtIQoSyaELjACjZaJbgYpx4RByzKoUD/xKeFNQ066p7GgmzXQ3m0UaIMgX20wQGS2qmGNgf/AKrTxhGJsgZGiWKo6kACUYEDwaqe+qoC8QEDYYkcMR/R0BEa8Y8FEQntCKtPcQgsoALlwCDVwCCkYqwBghLGmiDm0gMqwAISUB3uckW+KmnVShIimhKK6KkKoABs0BuTcBkGYR8DUSAIESIsYhD5Ya4LERnloALOJhCHIBCC5mfXmjF6lBTZeq81URUbwQSz4AaYsKwCURFCASgzUSDVkDj0ShNFsAsGBZ/86p4nCqIE5ao3gRz3EyoIARzlUA5cEQt8EAiTcCAGYbKk4iIE4bHsOhCToCMAUA1j8SMo2IkB/1ALN1sMxRAJUKmzPquzRRIJxRAAhPB2QsEATqIdUTIQFRcpWGSpikJLVHk90QAI6ngQIWIgD8ACVAAM81MOD7AwQSG2NfEGH0AAPICppqG2EyspJ7GvQSEm/1CxZiIB25oTA5AhILdalcMR1BULnSAvJEFdaQK2MVI5IYKwMDEnBzEWjccxhda2IxGVkksSs9FKApEIzhaUhPAPYSAEzzAzIqEMnuIpB0G2ChErlEMFXEEqBEEZl1RdrlIOI0A5/0AFhxMvlDEFxpALwGBSWSu2ymEcYwEOELFAdPQNa+AQdpCSlUsTegpbz3s9kvQPIfMPI6ACOaAGKjAFmaIGfP/QGAZxLaLCKQLhvbGQOsZAuxsrEFSABv3zNIVQCE5QK/FyU2hALulCBerzO/niv/9QBWjwD0MgCX1gC5LgNdH1D9A2BcREvpRRAtfyNe6QP7fqE7xkEyFBqYKBsdNrFKAZHhLiaAaRA6Dibe7iGHyQNgahAlXweTAcDM+wagYxDwixCTRkBzwQCD2QK7dbwO3DNQJBBmRgZbyDEDzgDpJgCJLjNAPBB9ZSIktEPF0bCBUqEHRLQXtACTvFEbQTqB+sF3mLPc3HC/NDLpYQBMBAUt1wC1nTCQAUPF8jENz7D7HwDOAgsbITxAThQ2w0OqewAOL2QwMBxgshO/a5AAn/NgY28A+KUMAA9A9q/A8pkAH/o0RdKwljYAdrULHfIIpV4kGLF8YGwbfGkrQbAcoF4SV7MQuu3AIjhElr7D4khRBDwL8FPBAFdDTYWwXkQBOFRagCYcgd0QSKgD4mRAUZYMmSw07Y+wy6sEAVew/ZsANaQMrYLKkgdDjDYzwn9EkptBCSgwzhoAu4MKhZoka4wAPpDBOPWxLnw7/ObBCSA0dnEM0LJBAhrBCcClTZTEEh075M4ZjjcapV0gIcMD0cEEmXVLtgZAjBQAWapBDzPEXONQWxoAPptUCaWBIu4M/Te5X15V4MQbCGhBOycBO2tEgs/Uiz4AfGZDYybQjp/7MQnnQQN41CCFRuMGHIQRoUnTADU8AChJAKDfANtHAHTIBtrkTKJ1FFC3HBVHUP17AXr3QtKbOpg8YGuVACCsVQoAJG5/M0ZE3JoiQOkiAEp/AO1tScBdGEL2FNA/FR9EAPZiAOJFXLM2EJaFAt8OoGbsBST3ABTMAEJaACAaCrkUJiwIKOQMFeTVERKtsRpvwPXbwQnOpTHLwQEccxDpHFTZILG+bVGBQMvJABE6VcByEOfEkPmXCeU2QAbzRCJUAJvNAKLMUCAqAK6eUP5PB52yer27edQ2U9FUQSHjRj/4wQnCoQHKANvMAHTEBMxDQDwWAAq+AE8umeoxQEZv+jBjOgBiWQC8+ADgv0AxRAWZGl3hNQ1GGFCCDwAgjgA8PgA/lKVcRmFCSNEgXwWhYgW3WRCJJiHDMRGgshd1zgYybyD/hSfx1DYB2h2hK1Ecj1viMUT93bWJWQCL9GDuilC7UAAp31WaDlA6H1XYsRC7+Qz2zrKPOqF0AwlT+x2QlRHc5mQTXRNwjRcNqDPRwgExaQC4nAB7zACN6WEIP8qhDWTDmdvyMENicF3pc0A16tYcZELpgjBODwDQ1AR/mspxcKS3f7ErRqEyDNEJ1d2UbxH9rBtxjUYg3FEJp3COByBXY1doLxCf8gZQWRZKSg50DhZUkh4QRBfGFmCa3/EAzWfcLlYlQM0WZd8Q+VMOmUsOE4Ra0UouZ+Y9JFYQFFkHQ7YAzDxDRPMWrY4Aw++g+f0A3fUFjYUGrf0GQxgA3+AG5BIej/kHI54WU0jOsGkWr7YABjFgx8ILJhVi6G0Aq58AS50Owm0ne0NgNEHg8pAV99dhSaihQGKxhnXhDK9g/KpuN7MXEJ4cEpcR0FUR28UDLdtt0cGRT+oBClViXoZm40bBBahhJdRm/4Bmv8lr9oMAPZFWYl8w+5UOkCAdkUcrVOAbV+M7MAcj0hOHk8QRAtkALisAqNjOf/gOcO7hOTFqmAA4UpcQQn9w9SiHMqT28sX3rbkAGFkAHb/1BvR5AH8TB/tFMjOp+sBAEhoxwUs5Xf2mGJZX4QnU0TVTcOiWd9FhAyT+AHWdd14GgQRch6JPcPspTkKBHvKNGRR3HyJ08TCSgQY0gHZ/gPMbd7MLdy/HAFbb+DyLANVQAMy/4EDyILhkd0pXB4ooADFrB0mi5XvbrcP7ELIKB50iFwyTd6GQBvNycPhZAHV+DuL9GRWakQl78QHB8UvYd7+1eAHjH2ChH2/6CFELCD/LANzLAKs2B3eYd3IBALTzD7GPcPXdAFr6BsS78RdiUQPy9F0TAbEosSAs0Ug+8xuvUP1hYIsQD1PtYKNN34pcfyMxf5X0oem58UbiiGAP9oe5+zf9RHfT5h+sDHjMhw/vzAC5bQ7LmQApwg/oS/EfZbreT+D7L6DzAoDmjGBQ0IENtWQYDQpg0yZP8S/mPIcNuVf04ibmPoBEKyhhk1buTY0ePHjUlAduwG8coVCMgKMoTQsWXLkQ170YHyL1+ehiQY6swZ0yMohvyODOEyRJyxN2963HGTy4WCBArUiWCozgPDNwzx+OTa1etXsGHFhqVAaCzIXWc1BlLLMUDDSJE8EuiI4p9dhhRcVTjXrK9GeisGeVzQFdbGGhlXZEzMcbDGk0cYSv4npvJCjTAZJgS1KtAuX8+GrAKVZxUJzR5xjsTZKyMJ2KVXVTnzAkT/ANy5c5P7QICAOAJyfBM6c8kXHl8CfF36lzbKMzltpU+nXp1jHECNNL4dich6R7nW/lkT/928eWqw9Jyr8E+YMHrrhOkRtvjfY6/0Gp77obFZzB/60iMJ+wZxpSFf/qkCixu2MW0VhTJKKLXUMuoMg0BQOEMJJTLkTiMMPvgnjLQYKuYfX+jKCAGO2GIIBOtc9OpEtUBAgblazmNIRh11FKJHtWhsSwcgQfqFFoZ+yZGjG1ypQY/FanBGo/YaWmej9s7x76wpN9JSP4a6sY+GfwRpiByNDmQonBFpqKWWE2mM858x/iFSCTsbIvOfOhjaojq7hCxyUARN5ApJQr1a/6OhaKY7AdFfEt0IkGsYiuOfNLqiJZt/VPknm18irU4XhuBgKA1TGboGEkgYOkEjTxkiUwdENHElnCQyEca8KqtLYtcrG9Jhzx8b+rMjMwFpiNONXv3HWUlHQuKfwv6RIlquvOs0m1i7UkWVVDRCx6dTGuIh0QZGWvSrVrHNdKxYw+VKE48yTbUrOKRJgxVqwXDij4a6ySiTf0SSbtfprgxWGPmCZQjhLaSQYlqO6M2I4obGzQidSGOA1TxtGYpA1YaU1ejaf9r1iWCGLJ7O5Y0i+JYbcTtCmSFuUgHnH1JJ/QjRjuB4hF+G+GXFn4/WNS/djoie7r+M+uvvH5rlbf9Imn/u/UfppqVhxWl0N+L6HxsYsqUhM3BtLInGMkoiHEYw6gUMM7rZZJOHG0oC75EW5ioJtg0OSXDXeunFBle6IfCfCqD+6tKGwpV351ZbPXeja1ShmaEuuQIb266a6fXmmHb+SGU4cEnjkX8+b/110IvE+p8iYh90EdujFSD3s8oYqVpJo2NoAt6LN/54kNa41BvkM7qq+SJ3N35s6L1ioHrssyc03WkykoAhGLQXf/yvmP7HfPLTV3999tsPqwOG4G/oEBTWWMOOUvFagoWM8GqoxI0owH0DJCDyyuEV6RVwfU+In3mI0BFKxKIHFtgBAADwj2owZBJemUQG/7H/wX8owwI9cIMfOMGQD2VkCUAqgUaUkb0JcECB7DvgB//BvBm2RQbZUxFXBOiRQzTkhQ0phxcyWA0vNCSJbalhQzxYDhXMgCEjSFQJZFCGFeZwOvcgWZFaZYF/ROEfF9DiSFgHFjdsZHZlZAj6vhOVOWiDFyooxwZBqJEkLtEndbQhV4bokSmwIIiJKEAu3FAANiZSLaLiyisYogEFutEr4WvI5hQpHS1kRIBxFIcFkviAkSyxiP8AQDXu2BEvNLE6HZzCEwoQxH+YIiOosA4OL1lGRxIKcue7ZS81skNoDKAHf+xKDY14StARMwoDqA4TMoKHXaTQl9PMiAv+EQpq/5KPGg35oVoeiMjtaKQEsVABQ5bBEFWGJY/pZAgxB5XA72wlew/MZnWwWU+G1GN83TyP9L7wD/6B0iPG/Mcxy3HOgSaxgxc8pTs94gVlHIOgGznnMf6B0IsO0aINAUAaT/gPCowFCDHhwvr4h88BnhGlGZnD+3xywYyw86AX/ccDyjECQxjiH3yI6UcwuhGBdqSI1SglAARw1Nz4QjcBKEYkapGNYjQiG3EARxx0kYar6gIOa2gAOMzCkHKBJAZR2GFGKOmRkjaEeOkDYz0f+IKVxtUntBBAD6g4UBc+YAQ8pUIwdjDRggLpheV4wBB/+o8mloOwSvQgKf8RCDncoP+Xi2DAR+UKEnqKKHtvkab5JHnZIk0hhEREbDn4YAkqjEC0H3FoW144WOpYAAu/+GwBZSlL0N6SejqSZkO4+A3rZBKmPfKDHzKii2ew5bU+mcIU+NCJWKx2LOwc7XITK0TsdqS1HAHhLmqhtRleL7fU3K10hssQeN7ya1G460hHItAplGMGrRiBYjUi3ZjANL7LZYh7XYjYf8R3BHclLXyDCsqgMgSUevxHKmpbXvHhDp9tbZ6najte5EUgBuQIBBjVkMlMxiS+OcgBQ/C7Eeo+QLTlmMJd78rfEJaDBSMIajl2EAxDoKETOq1pfH0ci1yoVsU+eQMN4ODZrWF4I/j/OF4DWvUCMPZAyVNOMkeY2ZAOdIAQxlBDidXwjy//I8QcCaoyVktdFk8hug1RQzD4UN9AUBEN/zAEMAiskWAE+AHVqEaLdVqFf6RAEv8YAY5n0FwqpmAIVQjGifvbUwxG4btrgAMc7AAOXyygMOClclho2WlQW6es+9AI8fxQhVzw9B8zyAEfcjCFMWfkwKNtJ0emkAtGN3cKcw7GCObckCFIog9NeEZDEtzoFucZ2P8Y9D+uIAkqGKLXdR5CE/4giSqo9r6OmMIQh3jAKVzQgv/YQSACQSr8nacUt5QfR1oaaniLhWs8zcU/ysmQL5eYIfdu8Zsz4uiGOOIfAk9w/4CrcItbPMMYUzAGj/9BhY3cYtjGGAkVDDCEWzTkD4pQBLMV9PB/NKEhkrAzrKdoiBQcmuA1ZQjFGZLnYJDDdP/oHvlmoREJHy8B8WbfGXc5vko0pAWUILS9wawRXizaRWpgOlBHgGtjqHYKKhatOBrSBCo0Idgiz0jG+/CPPiwgBmeg8RSkyJAqSCLYGQ9YDNw+7H8YAOKKODjbx3ALcQw4GEGgQgqAsepAiHYEnZjBCNQg7X8Eowk0UBqEy0jGr1CjXBdm486pnC7llWeAfiC1vxkSi7I9tgqiDbOJNfL0JiB80HRgyBUo0hDXcwQDDMGGHXiwANUCwwAhlzhDvv9eJ45AgCcZYRPZ0EQFiG8DGBBP/BRunItoo6HXU4iClH8RA13wwA7ApeYeGtLCkYgia/+wB8/Nbzxe5KIVlJDiaXMxBBysJRjMD0KvNaKCZ6CpG5lYgUTi3/qOUKl/sANWOAUe0IUFEJgxqBbbswOf6YoxGAMyKASuezbkC4IZCIZO4DuLy4AgCIINfLl/cId0Oz8TPItYO8GRYIBZmIVcyClL4AUD4IV/EIcUCDRgKIRC0AhAa4hoowLP+7I704gHbIgSJMIBLBqGwJ8i5Ioi1LCyUbvlg7ggeDhgyIBA+4cMMABDGAFfWIN7aIBF0ad7kAuO+CcVBBIC8z4CSpf/kMmdNPKKJmyekpoFPxiBGbACQrME3bOEfwiCv/s7jbhBYMuCITAALlS2MPu6hpjDaNE+j2EIRThEi3s4A9gGA+C73fuHORuBQEiDb2AazMsR/9II5khDHSkBZxqjaGmh2kHFaJkAFuSFAVODGegEAxDEf9DFjhiCjhsChmiCEMi4W2iCJrABkasC4JsOVsAFoxmLLLgCvws0Q6SCD/zAjOg1YwCHMGQI7oNFcGSj9GoeGWJBS7CCAWuFIMhFjuBFjpAEZKgCjzkXsTtAHmAFXSAVfnHEsODHmDAASciAbcBCi7vGjkgtY6ifBlhI9MmB0osJNvgHNuAEDrAskGiH/3AcH4IRr4ycDhZMBDzEKUtgR7DgxZ75B2fEBZ5pRrVQyelgvj9kiE3UiCrcqRGIghNgyHRJFykTC9wxk4/ASIz8Bx+Aho7UoivyneYAncnjJUNhMPXhgFmghJAMBktIAUqYP0LkHZf0R0npwhEwBnTgKobsliwauJGwJjbIuR6JSIawSJQCo+/5CExgH/DDlrDyCGTKnuthAKmkysI7LUsYMJSbyY4wTJRCgxaLAl1ogDBsgFS4g+/Tw68olqPMiDUKi728zIZ4ReRhQ9zhAAagxcIDPzzshBQwgK1UMkEEhsIbgSr4hcdUBU9gAia4S87UCMfziN6iJsqLiXVjiP/gpA7mKIJ780zkmQUumIHCm4EleM1gQMSt3D3EbAhg+DurEwdxkARxMAocIIMhIIP46zjz+Du5i0mGqMmzMMxgUAMVCMvGTIVneIInkAEGys2z8ErzKwUHcIB/GM7puCAggCu4qp4wIAA+YM7mZIgZGMnV/AdgNEyAJAdIiIZ38Ac90AMw0Yi2GQtGsIF1yNCNoAczEIdNrEJ3VIu/m74RiAVyoIVnuIALeIILkAHPO8GhpA7tkKvyG4+OjMhDYM4yYE6GYAEHhdBlywgD2E4kOIVm0A896JENZYgprQEyMFGGSFHqCIIBswI1iIUWkFEZZYInKIEeEABl2U3yYUP//NwIDsCtN+2lsxqJb9SRVdyIIcgFBVVQOuOFFFC0G7y4d6wAEU0UWJhS0AHBWsTDFqiEPWiFC2CCEcCDsVxIlcSThgiDNrWOulQLyPMJtrwsLioeZuCFGRjSIS08q/zTIbjBB4U9J+gHMwi9RNmEkeGdThiwAcsBSuCFPbgAFhCAseQqSCCEAeiAFviHteIIMZKrHNUiNh0JU7itTRULNmCGVJuvPUVNRSsERjhBA+g1WxywC8gFEMgGOAjFYh0AP5iAdm3XAaAAB1uDE4CRK2MIqqhWfc0dSJoONpAhLtDTBGXOWBCHfOWIwojE3JrJQP1DNOjSEXjPDyAHOPgF/wKYAIx91wnoACzghoX8BRR4AS4YBg1oB4w8gH/IUS4guvXZgJF41oxoqyEyrvXBzX19JOn4V4rkglZohRkwBhpMko2YkpFR2Pa5nPMARjrrNcMzvBxggVzghVlogQmgWj/AAmkQQ1XAA5ElWZM9ALAF23YQBQZIhE5xyvFxWbCgMIZI1h4pxbO4gJ4Ex+HyAi84r7ZQSpyrLC7ghfSLBUvQhpBSsj9tiK18VY7AwobIxMJTA6nTtebqAXOjgQ4LhJEVBQ3QgAPwgc09AA1wAC5IhFjwhQaYBobMTbi9HYbALa8oK7WAh4wwgVL7hzjFFqjkCJgdCb3NiOthAy6QIP9xeAI+oAiM+QijzR7SGQvFbYsbtIRgMIZAUAPIbbEpYLoBy0OCBbJeTQReOIQz0AWy1MkGqNP06VfqwFuvSF3zYF1TcEtsgd2PkKF/4MhLYkEGSKseOIRciAWIQNh/UNjjnY6iZaPlHYlrDAI0kL5gyEA83NMZSNAELYMWjYUqUIJf2KoGiADh8YlRLSN5Uh+47IhWYIigi1nQ2YF/yIrsQeGwsIBAyIVUG4IrWMCMINoeCYE/ABgjYIRPyAjXyAhS+IQe7mFSkJQCto6ZFNRBHAJeAMIFFlLmpKJD6E5tiAkYYVsMu7dECeGPACeG2AEQYOFOE+NYWNvHIgReoOD/VSADakGeT+iFICYFOC7ifyDiS1LNhjhihthBxbUEQ8jAKDaEFqjihpClcFkDXfCFQNiBHVABPtgDSsgFSqiEQV6pAhUfL9YIGKnWHcCEWIjkWGAG43mEbxAYhjACRYiBd7hQe3gEZyg+MPiEPuCBR0CaMhoCPU7cf9gHXuiExHvgGeAFZmAGLvjdwFtkRrYAFXiCSqCEC6AEouMC2T0LtT0/TljWmwWLHVBhSc4FSyABCrBMkIiABbjVjsAGr0Aaf7iHbgCDhrCFGOA+dGYIf8AFbMAFf3iHf8jL45GHmDhcjsiChthBj8gAXl61PHuufXDenQLmBC2BGYDo+ZqF/3TgCPHziWpOFAAan7VcSy4mlC44nt6Mli9gW+OEgRYIWidYxo8w5+mwZW8k5dpDHsrgCstwiH8oBIHWCGDMZZ8g6H+QhyyQhwyQB0vwWemLhWDYh4V+YD5YP1525ozwAVREX9vBLcriiP7sT+yZhI3yCMuzjg9uiCfYg6FrgVUovjaGHpiOlpqu6Y9og3+Q63+gDLiWjprOgiPQa3k4AnnYhhSwhAR+aj5ws17dhxYYOqMUBVHwgXHIZh35aLWAKQ8q41tCwzeQAAai0YW+gkJYRoopDOABHZfkHbnGjK646+84Atbea7/OgizQ6W3IgtnehxSwbdzOAN3ehm0Qgf94EIVcAgn6lRQs1lerjq2YuKciQcNyItMnGGReEIdvZYjiHe2OvOnzEAPtFoMj4G7ubm29hu2hHmp5QIg8iIeagCRRCIU7wIQ3cO/GMp7izh4JY5GY+FTr8E8lG4DogJEvAAB5AiNK8gM5ioUUwAngm5YqSV7kse6YYOOxoGvzIOibPm2W+AeYwIyFOG3LOAJkaG3WVolV2IfulAVRGIdS0IATdwBRQIBAcO+kiCv7BglO8Rns6IgZN4+0UgsVwdvjbgt9gx4WeIJ9yAUDyIC9hoDVUJ/O8SVkIAE6oINCGAIZXgXTAIU5oIM56IxtEAdgMAbo/Yw3AIFYeIJcuID/SuAAWWDxLhCF3+7PDR4JFslxBbrXrtBPr7Ds6ghpnxjHXtqFrCgRFfBbb96H8WZtMciCPLgCU84tuq6QjSCIs8BuCQk+EuCMdJiDVeDtYuYCQvgCEBhzUR/zMj/zRICGNRcFBxgHFv+HV6i3Tu2Ivsytn6MOPTceP88hEKgCLtDOF+QDGOQFeSDqXAiCFNiGvi4EKccbluaSrwjgkegV82iJ4cNw1PAKCY+J4eMJ4SMICFiFI8iApOOCfSjmXOgB59uBHgCyJ/CDOQhpPs8IyVTBRintsZjvaDkD9emWjkDh6Nhxj9idW+MF50UDlMsAnfbrI9DBK1hyvkGea3Fw/0kBhXwAin+AjWp3iY4wiLn+CtT4eG9fBX7gB6YmeGjuBBgWhyoQB05Y8ufBnk02Hk47i5689XBs1n8ggnZlCHHgAuMyBlQrCl7IKT6gAl4wdJ0WaqF2bcmoaYlfa9B5etuJcjrA+CUHioxvC0jXCdTw9jbgB4LfxaNfheBuiHzdaONBQx2Jc2xhi7nlzF1/oAGAhm0YAkvoeX5ghpFHBn748A8Xg76O7Yaw66B4vUsahYZAhlWQ62wfCxIABShgvdL4hyXPjODbiKz/iA/3u6PngkOIhUNyARFIgASAB9K3vK/airTAAxWGbIZ4+2lyueoY67GWA3GIjgHgAk5o1f8UOIK+TwjtroycJoNwyARNWAAkQP4F2IRp2QQzkIjmwQ+MmG6fYIQ86AUSGAiVaANJ94rM34go3wigoP6P+P5/AAVQoINVuAJxIIQXuJFdgKZdqD5jOIRQUICDvSaN2IqxBoh/AgcSLGjwIMKEChcybOjwIUSDvgTS2BXxIsaMBHtozEiAIB5fAS6h+GeM0MlwFCr8c4ZQWI0VHS/WmBkR2ao8zwI1WQUKFAQSQQVC0Egi4U8SeUj8zEOHzpVtQ8RVoVqlCoVnVQjI4eqVyIczIS/t8iXS164oAgm48CDCJty4CfHItemrkcBI/4oZBPEvkEC1BmnUPVhSL8EA/3z/XSKIotY/yIUnHzxT0uALghSobanQzCXBmIMoG5T5j96/JDUdUvOwCtm/QrAF8vs3W8y/2v/aECzKG1QhEGgtEhK3as7SPAWPZswDik6eeArEJfT2L1KkAAHOEKLwgcD3D/+w/BPgy3zjxnjOOFRM+j38wnEG8i3GNy4WcgtxNEQMSGAxiCF0QnwFFuSXQBTc8A81wrAkkGgDjSYQNdTMpIdnArl0zkGg/aMHPTWZJpArnFm2yxmFrLLKEcgcIVAbvBEko0BHQdAGBLCBsk0ggaDA3l8DTRQFAeLggEMh21zBiRND4CAOVRQQcoMHS/7D30AeDPSCXyiUZB1ieHWU/1l7k11mIJp13YcQYZGhqZc1/1wDCC15pRmRgKRRs4IwzXj2YDNJrOCKgxUYSg89K8BSkGkrZPIhoAn9EJEzFeixwiAjNkYQBhT8kxMJRyEzW0MQ+JTHEOT8iAJhbSI00WIDVbEgQgTUseWdaCJoYCBA5vorfGIiZF02//3DDUZKFHbNP3EOZGxCqhQk2UGu0GNoM5m4UkMz/zy4ULcaGsThReQmtEI3FYQg0CWuEiQOrf/YcIMN4pBBAQa3SDLENkpescq/2xRyJAFVPKOqu/+EoTBBCSvkCrARE1TfXr809EudEsdHCyICleSwxgXF+V8aGMEacscPuWJGauEitP/OQDAL9CCH5grkckc2/xPTg54KJMg/QANtEMSefnRCLZAp7aYvv9BAwxj/6PDPAgQJUeCaDtFAbUZch/w1RnCQJi2aGR/033wQ0bJ2MRgbKDZBZBMESUInECbEyiOC3VBNwhRk8UBXC/HoQhQLZLbXeyskRcoKNfGPp55icFDWcYF8Ed0YEUjaGv90HrYdEKUCLCCAxKFLR9moks2vuqRdUBysIItOnXZLsQLLAyVBEMx+o/ktQ4Y6GPMmMqmyABICJf8P4ZPLtMU/GGgiJzr/kH39YIoXpIMU/2z+0GoGmX3RCtAPRgMtckccQQRwfe55Qg0UJP9M0ggkxfcGIqv/S8kQqa/9QODAijRk4goiCEf4BNKNwviOMsJYxwOJJoTuTU0h0zuIswZSvYFY7ARr08gWhiYXAuUvIVMTGvMIZxOgXVAh/4vY6ARSQgBeJAY0hA8c4IaRaazBDuH4xx8I8kOIyIyGwtidQAZhBldsQRPtI1D3/rE8hwDihQYCnBVvqBFk/WN0qYjhQb7HDTAapGPts95CTiGQzBVEjQZ5n4GiQRA5FiaK/zgjGTWiQ4HMDlj0U0gQB2KDfgyiBt1IIPMG0g3VJGET/3DkPyB4JwiuIwlFPEg3wsGIZDghHCtAzT8mZceqVe0hrCjIKfPIRrjwQIuTiQM6Xje3uaFO/yBpsMMeZ9nFXR7kc7gYyC//gYt3hO6N06CM/JIZFzlGI5gEmRQkJvUPVvDgFP6YJkKiEbpo6LABfyzI5x5Bx4TgAhfjfM8a1tCAbjjhIE4YRDcWKBAkFiQJNmBEL0jRi3/s8x/scIIiFKHI1OyugbxLgkEdIqhtHSQJZmCEQPaZj3/0IxxmWEENBJVIjKTtlKxA3SnnQ8ZWDgR18+FiQ0KHOmc2xI2Ks2NCZEmQ9l1Tmi4diB2O6Ur42G+npHGBTzNCl6AStahGPapDBIDUhyxCIE1d6kPgICwAfhOnS52AQCaAVahydSAyNVARivAPsRbEOl0dyCKeetaURkKpa/+lYRQZ8Na50rWuUM0TDauaEbPata9+hQtZ/yrYwRK2sIL9Y2D/AQPDMjYuem0sZCNrEzLdQbIPQYVNVCAQFWj2H1+NBF68ORCfEWQOA3GPZVOr2tUOFgVwSEMadIEOGgSisiwYgUEAE5iBoABwrP2t9uQK3OEaBLMM6cA/DiEQQqgFBCCoBgAOUo2DTGIg0Z2uBf7BgliIgwtZ+gdqf5Vdg7j1hlslbnweUBi8eEMveEWvRp7QEQUoJBH/KEAsVKCM6v5jugKZLn81Ul3//iMWueiBADCRg39IAFgl+MeC/xHdf/QPvh15nEM6uzcvDFcG//AwDZGbEdMKJAEDES7/QVRQDunGZxLVBUIPSlCCBS/YCgZ6MEEm/FsdwtEgai2MBGJRGARk5BgRCa+FaWhig3ChAIfI7z9cbOQCcVggHF5xlf+hDA2nqQwlKANByqvax85kcg8ZL9iWcdSeWta+F6HvP+irAAVwwg8sWLGVC5Ll//5jyixmCIFXjGeEeGEELPiHfAUiX/EkudGQrexAKuzogsA5zpwgQhEIvBAvqDnACiGwn/lcjUlkec8FwfMkdjCCXCR3IAgwBVAnLWu7HsINuJp1QTA7520QwQJqNrWe/1FlDuv40/8YNEHKMYnpKhvZCeEwhyehhlzkogACYQOus21XCZAp25z4lAK0/9FrDqvZ2QZR8zI4LRABTBjYUSbIMvirZoK4G9Au3kEsrE2aHABBIABIHFFBrG3KFHvgaVqwDEyhAGj4QQIrVq9D0i1sL/DXxQqZ90AIrOmZSJsXbHCBKd4zVKS+gA8GPzldrcCEWXAhEBs390JWfAx1G1sg8ba5pwndEAALBLcE+XFGypADsv4b5UZfbSgM9N4FX0AF/IW4Qqq88XRv/CBeqLrOMbJinr+B1QIJOVze8A+6FCOXRz97YUORdHNopBL3bTVDpoBbn3sB5gWZxMyFHeqBzFzNeY9IuesueIzXuyGeGAIbgI52wiY9spKmYSgqDRciIESpmBjBBQoC9f9k07sanK53OTi9bABEFxP/wLjdT696m9e9IWqe7qj9LZDqvsEP346PHBave8GynVcPEfSxyzGFcijb3eXuc5UJP5DC/3fZnzd9NY4x3euSnvQSrj4A2K3U6ArAAtQJOkS8e9TM72r3cnmvZSV/ERFfBPgGUe8DvDCFGQTjH6xm9kHwvIzQIyT17162hAmAAGiHdkRCMTRCNsSBAroOA8bW6ZxObL1WGsQBDcjBIngAaV0Ejs1V5jla45nf11AeQxzaQCAbxiXbDBgCFeTCDJQD1tWFso3aqAGA9E0C9pEeJpCe9pUHeKFWADTCf8BBHJyBONweRIDZQxAZV7GZZW3/wA2hHwj+w3/sgECs2BQgxAkKnyEYgiXwwRXyH5rMW+htnc0JWuudHiZ0GuzZoFsJwB0oIXAxAWt9gZgpDnYwxFdNxuP9lU71gG5pHiBWoRp0giXkwhXSG5qoFxhmhKdhwkf01QBkm3Ipl0CMHABB4UF029EBQg9wxEEoQ0LIXSEGw/Bl2Qmml/thhKYJgCcQwhnRFRz+g+IRl5sNxKZA1TW8gBssVhQCork9wBTEgiUEg88RxOYlxClqRDnsn1wAQCDYUF0xgFyBHYr1YpqEV4/BB5INxB9FQsF1hCMIxBfsYV34wT+Y4z8Ihi4EgidCBDDyASXMwCFehKlBXDk8/wDw+V9DHKPmDZrFAcD40FU1WmNkbaNBfCNS2c8JeIIK8KNCKAMwjkAnjMA8RgSwgWI+atmxYQTUOWRCAIAvmB1BjiR8DKBCiMneZUQ4GkgkgtMZ4JYW/MNKxh0w2p8aCIRHxpzs4eMDYORBdOQ/QBw+ntpA9BtCfGEy7kIenpVcDSRJLsT7SNNckVlH5CRloCMhpIIqPMM8zmRCgOIU4OMSeGHq+V/dLQNYqkBYOiT8DYRQTgEfGMJGbp7wbR4oCsRdHsQuoEM2/gP9kONT0lVfBmZG6IAxUGFMCoRXJoRYzkBCDJqzpaLw1d9N5qVBXCHUCV8roAEVOKZGloMyhP+lz/XkQFgmTkaZkb3BL4gkYdpEBdGQjlHlU1JlBlFYBHhCIFyhUQ7EYhZEWP7mRkZmCSpEOeDWFuIWUAqEGsyAClQZ8RnnP1DBRP7DFAzfsd0kH5Diiu2mzr2BL9TSQAxmaz4EGKHZeAaVTi0BQrQkETDXTRblPyTmUVLnAwBBTZpmFVJndW6kQNTf8I2AYwaDIeTCCNSkQByiGvDBDggaMKagQBgCMBDoP7QCRaraDBhAClRBbv5Dv+1mv9mjv4HAL3hTA6hTOn3OGpyJ0RnXP7DoeaYWa/5DS/5DC9jfCKjBTWqBGlQnd2pkQfRbWCrE8PWAPB7bFBjDPzjm/Mn/JRr8Q4Ti1nYG3wjEgjyWAwDsQCDIJUE8zi04JkVOQTBQgQFIAjB44QPI5zz2aJDUwi/UQtP8wy48Q9SYn/q9KGuRYAtMQI3+g562ABEQwG0B6AzglhrIpzEahH3qZv6NgDhQZEQawqD+oUBIQhXcwjNs5CGOgCGYHPEFQv0JBDAMgUDoyxAYwkR66j8YQCGAgSTEQoFqXpD6aN2pQCBMmAC+wRSQAzgIxMkUBgfIgp0GK7DAwUSUQCJUAiUkAi/8g31RAh/wAQuwgArcqBr026D25kP6KG+ahFZUoaYSRBVE5xBAABlIQhMYA54JH/39wwi0q0A0KRWkwCeAwT+Q/8E/KIIk/AMaBEP9jekt6AuBtqV+VmtQguJd3qiEid0U9MhElChSMUDIzaLEKMAcuKiwNtY00MChMUEltAJBHGIO3GSOviduVeRC1KeWHeMIVIF+UOR7hqu+psA/XIFA9EETVMFhDkRFwmt0SgIZ3MI/NEG+KgIZGICsAIMkAK2+VMGXqpfcOSuebV7JsituPcMuoOhRNdVTOaWBYNWeGsSSXSxk0cCDPZjbPcF7DkTaFgQfFKNCPIAjYCu7PsMt9EG4zh8VgKqohkAT2MA/9AHg3kIwLKhAmNw/wGzPJm0fEMQY9MEfZKhA+OtAUOqXrtgM8AIvGMN+BiXxJSlBBP/CM5TSUkkj2JxXroWt2ELWEmzgQHBZQhii2hoqh0KYyf2mI/zmFIQr4GpomApEIA0E0NbsGHDlsTno4TrpPyRtQSyAM4zBLVSB0QLDqBKEJFDBCKjaPxiC0f4DKYZlgs4AFZpc/QVDFfAl/JxvUXFtQyRa6iLVfEyVUbmZyTaM5k4BEKjAjl5mLBBCFeTC4E7BDkyBXNLBP+QBKcSGqBLELazLuozCAvAAOLiDWoKpvlaBqP4B4NZsN8RADIDDAozB44xpAg9ECPzCLQADv0anzPbnfqZgK8jdFgaDOARCydwD+hrWHmyWKU1GPbRvRCxlUJljC3BBPH6s1/3DpQ7/BB94pnzGZCwYTPJeATIUAh3EA0TwQOjYgR1EjdxRgTgMwR/ULUPkwxUoh0BMlEA4wQJggDhQgRsbwBDkrSF076p1wkQGg4HFglKKJ2Ed8UNIg2z6MHwEclFxAQvyAQvilmNuQjH1XJgSI0H0Wzn0QLg+QxN8wkWMgR3gghbbwQIEgjFUQRMArjxpCDYoBHMYhA2cMBUAQwYMAaX+QycMrqbmbX/uABXmLwr0yBh8TuW4kukKsjALhPhlVYEBaM/NABWM8D9QRyDwARWo4KAqJnX+hdW6Qzi003IkROfQES7AQQxowi+Awyj87SiMATSi8kHwwA/9gr0MBAkMQRUE/wH3amouRDOGVgH97XOQBEKMDjNABxWKcUELtEAuUIIiB0EQ5G0hEIJBSKdATOc/VKsaOAIoowA4oM4YVIG9CoQ8I4RK/UPofDMPLADhgGcjPwS9LsAChAMGLC47DEGG5i0aoMFCL3QKGEA0Z28VoIEkzGliBHRgoqNgedchLDEaUAIwBAEwWEL0FkJB5EKTynJ0GkIxXuEVYjROAaZUFkQxsYIdfJRVCURKM0QMtBIPbMICxMAP/UEcu7G+LnS8ZoAbiykvzDAc0E8gR9gNcQBj8dVB5LBGmMCvVBUVfo2tzYTAgQ0DcIF37UMGyEMG/MMQyINAZEAGpADNCgTfxv9xQaABpPqcI7ynRRjEP6eJ2PhtE7y1QNhyCmTBP2D2sv5FLYhWQQTAKSbmFwyzh8khXDiAxqiC6/5KMGsEx/zDOWmMd/ECC+Dogy61QZBCEAXv8QpECgzBQqOBz13hp2pEWcvFKQlEE6w2FdBzdAJDCtB13pY3Fcjd1epVQN7kcAs1XBB2Q7DuXM1o6vxDQH7NLHTADKgBbkHzUktvQRTCZmMYqIZqqEqCAfivzwUDOSyu9uzq5MaxeQdBZuu0eWcvuwaCLtj2QPS3IOMVCeYKfgPAFxgkYbmHJQqEJmoMis1CItxou5a3gTtphxtEFUiCg+f4uuwLlPivMQRDacf/hS7oAivgglhjRO7si5j+w2tz+I5b7wgEQiqIVg8PhOnR90AklsSAgIqzuCBPwCwgtICPAI7v+EFUgczOhouQQRBR+Bh88M1SatR8d0a8D3hGBDv4UyHotAFkdnkbBGfWXyCMqDfBEZh7Odh8gdillje8uHnRuI3PgCUEgQHkuENYcCFIgjv8AzTGgC5kNA/EwCgggZ6HDUtphEynN4b/g0IXBE2PQBQsAIk6+lIR8nhiFRfMAoEKOKZruiUQBKcrhJNYjB3oQliHNZMzuZKv+q/QszzIQwqUN5sbOm6NARyoE683BAdgm0McgK5DxDdwoyA35SycuY3zgQFouvQe//tDLMAmTxPqhLS0A4tCuzEwiGm2F0QnMOczoAOJ0k/jyKRDiHu5k0Yt6JRAtBDaAbdGqDuwtzsvODVTx3tDRDlBkBRZ/xInczJcKPlM6LSsE4TJp6otR6est8IO9MB72za12NhDwBpGaMAwdITEEleXpwkfL0QZLMGhRTrYrIE3agzqQgQDrHsuNPeUYm4QBANTL0SH07OmTwbJa48hHCmIN0A9iBYkvAB+yy7YcEKsmcLOC5bp7fZunxUiHBoS8vWdFDdT/sPS7wOBWgGAWoIlTCQVLKu8y7qB/7tgsbf1gjINFHwD/I/cI4T6xodf/4MLpP1f6Vjjd1UZLHbEMP+hLQUl82kPL9r9ulOC0w87MXYCL2yvQhQ7ZbS69ljCoI6AEni7N/1COy7B5R+EWhkhSdYhQ/S8FkHaP+C3T4mVmuFnyGDVLDBD3u/9RFoB6m/6ydPzsa88QVi9X20vMaqBMagC7atCFHgYjq0tQkT+P4AdQB9DMt6QDPh2UYlVWPX1LCTXDOj9CCxxu0a/9OYt6wPEPwP/CBY0+C8IwoMLGTZ0+BBiRImdRkwxdsZOA420okj0+BFkSJEjRTY4eILkx0kpWZJk8q9Ex5YGu8yEWOQfTpszCxhkwOzQCCtCiVrpxCuFOIH/gP1T2rRpw4Q7I9opCO4gFYIDqUZFo0b/TSxBGhvQ6sGkBEyqa9m2Ldju4Rq3c+nWtXt3J4d/DDjwimVlxtChI9BYMmAgBdeCTSUVnKowCDDJwMRVYSoJWKGdughadWdQq1aCkdcCozICbCwUGlVFeSKDSZm0eGnTPlAbd+6dJv7BqwvEoE7dC/X+44LA75LAI5YIDWYpRdSIksVRoPAsBAYKK7ZvX7HCzEzOBMMVrCIOGGZgQRT/E91SeivUOYydaJAKRRQLKlSwGP4fwAAFtMs3vHASbkCD4lCFkFaUU26wfyg5bCmCpGuMKwqQ8Cead5rRQw+GhPnnD1tS6uOffsywIYR/anhxhRpWuGEI9tqC6p9OZphC/4URjCnmlzpiuSMWFkoYgSABElzyo3F8YBLKiK6JkkqPuPhngCcgnGGJf7qkJLEUGhqosSo0ieaRd845xy5FagCRIXpcIQOY9jySDs/FFgsCtSlmMAaFOy5gohUmYputyijhSpTRhlQxKJtGJeWEgURYmAFT5QjqhELEChKzoIEoECKaZs4JMcAabpDEEsi6YgpWNOZbIhc3LrjVULQsEAAQSX39dclGCJIL2CUvMGiRf9jg5dJMvZyhk6RA9ZShJpB4B0RUAZxRqX9aFUm6hnAMYgY1UBthD15uxVUGFXiVi9hi5WXrGN1aQLY4iF5yCI95o2SDCz4w5XIGJPmg9v+hFKz90KEaahtkoXDbIvdcNSip5IJWBmVCBTwAWQOONaLZggAiFiIAJX/dGkfAY1ZiqRWS9DIl34f2VfmjXv/jopWBMbXin4OR2qqhIZoQphl6RsSZpSCCMResVijRmIkLcvB4DY3g+KWWf7z5p2uCpmSaKpbJnokNkp44myGT4gCQmVwwLQNTJGeALrF/QD3IgCGqyAQ8atgmic8RchCKD0ooqVoCrDVKpQo5/JjcjwH8MCjewTW36ViPTGGj5s0/MmlAZngRmG4u/7kbKTGj8vQKg8IZBcAKDtpCNwOCkI+oJSjZ44Iedokj6/sI6cCPDlqYvIOGcFjoSdEXYtn/bKb9I2iPkExJdiQZpBdQryHkTh1TCVM4/5/GvmfLAD4qHqEVXoRPo/hUKOjA8gk60H8CQiBpYA21AIFM1lfAhWTvIwwoiCkMeJfqsaQ4bJhFIgZ2JEx1whJD2EbsChKDBraEFxSDGvyMEYA0PI4CftBfC/a3P0KkAoACtMA/nlTDg5Tigzlsi/d0iBs2+GEGAhNYwYKxQYP8Yn3qs4k4DGAJWY0AilMYgRvIoREeEECFWZyACu/AihiCQAUIkIUGNPCPMh5EgT00yA4ayAk1+kovDMiFwEqgnFisQikedIge3xgRXiDkaRVjQSyegQIsbhGRyPOEFxugChBYgAvD/yDjASjpgwO04wAOYEDn1IiJf3iyj6EcSfSoQqll9QxThjiIFBjiwR/gbDx0SQwaCva+WPiBF1xowQR26YcWeEIaAATELiyAAElqgJLJ1EA7ZLFJY6BjcHBZVEQIWKzriZI2PjjjP3DokRkgiiAMjCMvdCQwefxjAa1kGh/dYieCJKYTwYCiuaaghin04AmT2+Ivg7kGQOABBJHUwDiSaUlkOoALlSBE2EjXqLQ9ZJoPUQbOZojNlnghItsUSQnScq+9HCQRlogFH3JxhSb8IwIoZUhK37g3kQzEAE+UIlimUNMRzIASd6BFGuLQiEsAgAtj1IAPLGlQDbyCAZWIRf8tyAIsNzikjA9kCBvvApwktaQnBHnBPyqqmwmQDaMQkepHwOkTLrjBL3zohElVatFP6Y0kGTiIJQpW03o6YgoPKEc5prCDQIwgFrHgwhzSIQsfDMMH8/CBKDRggoQ+gakAbOo/Gvqr2/zjsgJahlWp0oOuPoSBd7ncvMK6EHg4YCR8OMgffWIcFuTiEE9oBQfTiRse+ANKLjWIbh8iV4IMwSCWoEggdjAFvNaUr/Wk5wgSl4shcEEb2gDFKrhQgKWSBbuVtSxmqbQM0RoktCPhLEtMwBveMOSrBYFBAWdBEC7cIRC5yEUJMnCFTSBxITGIADvdWjSHDIErTfxHLgz/UVfj9rWmYDkXYG56qZvGQr6FBEfxsFuPaUQDDtgEgLw2MBIEDuea3+PALK70jzucrqR/IAgrCZJSD+q3rbThwbyAy9uHUMEQtKzlTKEIRZ+VwGfM/cAtfJERsjSDAv+4wUdY0d9/jFc3ofvPeQ1S4oKwoBr/yLLorkTif4BgwLmIxRAgMIZ/sPggMaitTXD7jxkTJBX/iDM43vxmiPBgHQIago0lEpWEJMQwlrBEEDrRimDUbW5BvlQuCDGGxxmEDeF1CA0Iwkl5TfQuaRTQhxfyWbxQNVFvKIgEFsIxiLyhB4cQMz/IwBA004WPY7AFGP6g4oaA4R+fyLWuDwIG/1zPBbi+LY3EDpIYJ6LypjMgH0kJgYIBuNGNIslFQV5Byv4ioC4M0DREnnAsPqjhk6DODSgTtQNyG+RmEFFBLA4RiyrEbgG1ZSlBnBHjtnyC10awdUOMQBAj4Ds3wu4tW+QKXILwgheUMESyh/iPWPyRGR55g3A4LeUcerog2KYL6P7xAY9kVQUBEjeV2EjVaR+kSxCxQCDEQYkxi2BARuh3Q3hdECOQghS0yUAGDO4WYi8kCwU5p95SEM8gzuAfIwgGL7TxDxcoayHo2AVB3mCBEmCsElmvBBtwONYCAgHjUTq5k+1C1R30gBJy2wZBdICbXx9EEYr4R791rQhf4/+aFP+Wec3/wY5G6VaJP/+tRCyBSqTP4AlMNwgBaNAIdFzDF2/YwQ76Y6hu76ESHSaJ5p/+K+BA+VdmJztVPhuLRJB0QN8gCDaw8Ye3/wMbuMDGN2LQDbsb5BNjwMY/NiGpnkuk5wIniG/lKtwZBCNoSJ+FNtjABiKo4A3R30HVKc8CtBhKtdBIyQYk7SudhB1Ke1ibQTAx+dGvZYZvmEIuOjFgEhRkAa/GyyMIgot75Nkga/7HOx6BjU24PgSwwQ78QfbabHCGIOgaQvg2ZXUw5eEQLhemRsyKhAWQ5AkuhhIkRGpWIbNG4qF+JeSejDai7R+4hyS+QHpeZkC+4Av/3gAAVCDt+GDtPkMi5u0hHoH+DGL3cvAg6I//sMEW8s0WrMIg3oEgcBAbHsEAa2MBHaIJRUKunlCu9oEXCuzQ/qEVqFC1BIYghuibmgWn5mAYDEIDREFSog+Owukfuu/8BKT8QOkNAuGPkI8g9I8kcEEkjJD+vsEZ4o4g9m0hjNAICTBRjsAgnpAqMkAeLOHQ6JAS9oESMMULgUwS44cgzOayzLANWYIETRCblMQgSmtAQOAL2CgXEu4fVkGJHiIC6u0hdg8k6G/33qEBnCEEQqAb6g0PdfA/EBEijiAKF4LPRiILMqAY98GJji+IOgEZC8wLgwjhHEITGWXk/sO7/yKCDd2CE7hn2w4CteYFFf7BHGpjB1iAElqgFcSBgwpC/lrMGWyQLR4BDx/hHoyQaRKwNrKgGOWhGCkBDYKhZ4LhORCuFSIQFQfMyjBrHjaxIepFBQVkEdKGBBnivAoEWMYRN4pgkCiBFyrByuzQIFjqHV2xNngQQIIOHyMiJefCEA1RH/kxC+SBCjuBDw6ND/hAahCuBRSHINJmGllmGhmSSvRiG2kGIkzgFRLFC0DRIMIRL96gX/7heiqhBXJhFdBpxf6BJBkCJGnDJHNj6AwxIpDhH8jSLuRBLP9BH49AH2MyA1JAuGoSJ2egFY6CF/bhH6YrHV6hC/KgC/5SKP8bRS84QMq+MSQ2DC8egEmisiBagBfUcd9s58wEhP6+MkHEwCAw0yDEsg1oAyXZki3X0i3lYed4YdCEqxMMwRCkhj14YQgyABTo4BUIIDCvyoC2qiAQMzeckiAUgDYAQAK8hw8u4DGHQAQ+A81YqR11YwlVxizZIi3V8h+OADTRsi23QR8zYBuMURG5sxizYBvyIA9EQRSSUssI4twIQuNK8D/ADy+Y8nvcgI02DAAAID1xIxTq4j4lAJy0wRKuwAnQqSvvAhb/YRcLaOhYkjrRckHZEiazcx/BMzzjwQxFoZtcEBOq4Q22rDYfohsHpCYeAkHoIgeGo8QOgSEEIOT/+ICHVoEXSkoz4A83DJD+mnNwqNMtkEEsMZM6j4BBfRRIr3ODVuEVKJSxSkEUHCAUAmFDXbBDHyIhP9QtEtJXcgDcgEAUaeMFdPMgeKgDoOFFgYERrKUgJHMro+TFRCLnRuI5n5MuOhMZnrMzDwIZ+KENeJQsxeAI9LRHC+EItmFPV0EbQuEVyLMMNQBJHYATLOANMOENpu5JI2I9IUIGNEYkpDRSAQBSC6KiSuAJEiFuciEFSGAd04mV6s3FXDFN75ElkKEN3LQt2uAIIAAU3g8C/gEC2nQ6C0Is+WEb+HQb+IEfVmEbtuFFn4ALChVJE7UUHAABGFXURC1SGyKN/9LrqRwCzFSrLhJgScoKStaLDxDOEIyxEEDB71apIOARxkQJVjtzTqnCEGmVDvKBBEhgFaaLBCBgFfQVAvp1X/+1WMUhFnbAAvCp2wqAAwrVAcqzPB3gFQZg+jo0ABTEIQYgJLR1JyYgAUJ0Wp/l4QTNGLOALelgIc60Y0liJQmCLMlyFUhgCILBGLhgGzhhZrdBGxCAC4yBSV3wDQTgUS2ABS7gCSqhADZAFkohUUWhC1BLDjwJBRsivaQHB5aMIDxuIeCzLdbLLjiW7KaOMXdgBBLhRXmBNEXzCOig1TaxDW61Idi2LTTTIHIVFOaWEzgBATjhOLjgvaIPBKIv+v/wAGiFtgAKABpewQGQdGm5FiQw9WQL4g6CxlsFRFq/BwTwYOriEOE6gRJ27jtFVh+RIQ+aIJ0GFC/gkVGQoV9v9f124l3boDNvtV+voF/tdRXqVm97gGf9FiqB9gm6rRKgIR26wHC7YBqt1iGitnFHQmtzIwAiQYe+IAoIQdUs4SY5khcyQGap83w8FwLyoDyeFALeL19bYk8L4l0XYnX7FXXLkueGgBmoMBZGYPL8FgTwKRaeoAPmgC8BkyUsVpQyrC2uNXklolsKAgXOIHpzoQpO0RIQ7jVF6hTlQYL5kQQY4R/MTCivYG7/IXbC121Fgh8g4nVxdXzVN1f/gR//5IEXgKGBU4AKX1S+pu0U5yABXoFbDcIDkjcN2CIWoGRi75NRSO16eoAgRst/CQIFCGLqAEAApIgPLIESbtIQUkARPbcQhiAPApQlAJHe2EIKTJYubvU5SYAOQIGEwzc3Zhd1UxcChHXPTDMCrRfhxEEccGAIPEABzLMgNnVJJhdK4CUa2EIG1qsaT/ZpD8JiiaAHQKBy/0EAAGAHcgGKkS4YDCBk+RFIC0Ez0rZMW8J0ZyJlACQ2zfgK6pWDGeIqYTdHU5cfWJkffDQDEo4SLiDteAEBNE4OfAXMGoiIG1dYGoJLFyIKRC0KquAQeCERgoEPDAFMLjkmPbdH/yEP/y6YSuqNldouQN4vNsu4Xlc3JMjSXf8hnD8iddd2bXP1lcWBCiIwF7hgFfJAfwd4Lnqgl+X5IPxYHLggl7gAb/WZCxQnNQ2hgTnXLdtSZK1TOhtizUJZN/irVXeCDiK6m1NinCHCbdk2X13ZWzCIF/gBGkQA5ggC5nyTUTZ1l+35jcBMDsQhFKBBn+cY4a53CKjzlYP0QYOuJVty7SQCzVagdOEVnDszhD9YJGITCiRafBvCmz2CqBeCbdv4CMQBil34rD5gERJAARJABBLghnPzH/qFMdUoyVA6QA7ZkcGMCExGHGiWC9pZG1aBH+r0TvkUR88p6DRDM1oSLQuIdv/SNlchoKIfYh0ZwozzMqIJYpoZIqlBQpUJwlYJYl+3QRyGIJeIwBj6g904QQSymrNFID8JQlP7BWvJhjYlYqz/o57lOZgLIpedAgGKtTiFNVfn2iDWbgim9gYoIByaoDwKOEBgoSEER3BG4grEM1fBGbBx9ZRtwoxJFrGXmiFgFX0P4iqv0o3F5wx2oWffYN3u4BA0WwFIeiH65RJ8gSAmlqxFQiZ24RI8orSBJbWpQknCuiBoM5fFgRAIoQrseBuGALhidO22oRBuIBMWwBleid6++B+aYTmpIgkIArgdZidg9TnXERSuoBCuEnVRN3Ze96k9ArofoowT27GXm07/ISB2YudeRzkPtgEHmk0A8MByBeASLgEFLCAKXoAA3CgUPNshYvwfzBtndqEKPntecFOJvwc3PcEt0Ptk/sEyLoEG8AAFUOAZPkApirVYr2AFJJMh2IQe6IFJgPsgcpgh5AEzQ5ghXhcUquAZtgEUYnd8Q6KwI8KMSWBunTuiIzo252C6pmsV7jXQr4BYt2EA5IAAEJ0AXoC9d0EAfCHGA2AXXiAKooAAPMDIG4iPi6WrNj1K2nsnAoE2TnshJhbMUOAFDAkDpKAZ/gHBm6EV/0EPkmAFyHwhkEBAbJ1NVTbQA8EXWE6D91V2CWKwqaLOCX0OREAcCmkXIiEAnj0S/5z91wngEAjA2q+92XYhAPAgAHwhAC4hAJK40uXAzNObLUCdIKoJ3Vmi3LUYJNAdBSa3a+jbI7bqDKgEzMCMAFxhE0zlICqgAmpA1xeCdCFi4P8BuBN+ISRcImIUM8UA4sV5Id6VLEGhEALB0f/hGYZAg/9hzqc7xB2CxAuCjFcBB57hH3BTAJzd2aE9AAIhv6+92qug2cDdvL3d0yGC3s39IYrhH2qcIJTAICBVyP/DeX9+3f+hGGihSo6+JSjAFVwBCQ7cFX9AD2ABYvCCHtZhTf7BduihGwqC4RG+IAYht6ugTv8BUBdCDJABM+d0Toe6LPMSB3zBF6j8H+KQAP+GID9HnoNC/iDq3CDiIQ+u8h8C4dQNwnkXX+lRgBA6ruMIIcmw4OfZYmKFnud1RumDPGzuYlJzxmu+5msKovOlJ4kLghoooAJMxVT0QOAHIesZ4uA9ogbCfE0QnCBanSB+wB+aoQKSoBscBrh9miBc4QYwIBCSf4Ne+eHF4HwN4jlvdW2R4V5xAAV2AQVEPfkxX+OrYIPg+R8iOg/2fM//YQ7yABReQTy1eu00Dgc8IdX/4fQLQljq/yEefyYuofR5niAAIs2/f40a/StmcKDChQsRMXwIMaLEidYSPiz2r9bEjRw7evwI8ca/GzWaSflXIcmKgUlqqPzXzxXIh3r/ZjpTWKECvRoKYf1ztQXFvwCBCOHYtorfkW0D2/xzqhCZQggLISAjAYrTs0CBlPw7w3XgpTP/CP2jQKgKIQx1UFzyFSCuLyw4FNb9aHGm3oWX9k702tev4MGECyvsS+sfDcN6rTF+DHkjCAwKKeT8d25hM2ErXNHTWcPnyoU+H9KbePOhsx//WA90nbnCutD/VqzwOhALoWdVxIX6l+efVKhSB0otzhDZKlAiqgRCoQQ6nksBcCvEoLvOQF+1fP3zPlIiWYUghEY+D9K6RvQKve5iDz9AxMAa18M/+C/SP2uAHHvLr999MwkkoEKD5NRMbP8I48oKCGL2TzM50ZPE/0KD1FCDHjU189hNN2X2TyaDZDLQYih4ohAWFAyEwBXAkUCCiy4a99AqU61CxzaEoOBWYCleNJB9IjE0ZIFGbvSCQvYdySRhGJnX5EPWRBLgfgPlpVAchekQ5V4yCVOBFBX8U8OFHD40ZmapCaOhkWHi9E8dPi4UxkI3kHHDNk6EcsUqLi63CgmB2jgQKP+sIsIVIuCgRAC+zBlRLcVIuphEIvHYJZNcBplpp3tB6emRPFYKapfZJDaRK5rocU4NK/BUwYcSjclQmkYmceZQC9UhyEArQkQBBnE56gtXSgQyBrLQYSoUDbUs+ZB1glUaKpMYeYRqtdpuu5CWhZXaJP+q10Z0wxYrDFLhTLRG+E9qD6nZ7kcgPjRaJpQt2WuvEf262KTFXPuvow/RQK1EQnBU5ETQerQwtxPJ57BhBIL0H0MFh2qQRQZ5O9jF7KUy06b/1BmsGWbUAC+acKrG0bzsSiRFggu5e84K3SykScX/HKzJdRA1sRAtpypZjC+/QIkCeAwpoW/HDDU80cH/ZBuxYdlU/dAaa8ARGdVMXq0QIP8AIvZAHH80LpNpxOH1Cf+c9JBDpAoSxg2u8HTkuuqitOAK6wxU0xb/uD1QzwONNhHY+HXkNbcib4T4Q6pgHREkIKtygsedbg3HxIRppMrkRzYOyDULef6RY/+ogpH/QwIKhM41og/k9tkDub7YCVs0KExkLqPXkmwNCYYq1Y1TDvc/XKo+UQgKRb5QJFAXhuVeqVw+0C8gJX+e1l2jis4/tht5Ddlm+5VNNqpYo/hjBKbBtUJc6xJHKrIPFMFCusTNpSu99045iJwjJwCsDBK097aBIEFqEMmEvgCRvn9czSCqON62NKe8x9CieoxBR/gicwJIMSR/8FlDR0xowoXEbyaEOxIgQOYXElqDFmWbieEmwjXUQWR2aWDFP3SRhlQAwiERcAcOBBcxd20kJzUZCJhCBIl/IEF53PvHDUNkxbENpIZiQ8fsMnKC9ViwI3gbiDsKwz3TfQQDSJSc/2DKuBBnPQYcenHdP+womBRCpAEP4SNDUBhAiHxwIDrkCDrExjyO3LCAkUnDxOKwhRuYYQXpEtAUIyObdVWgd7bJ3OM6EjuIqFF7DmmhX9r4kRpGxG0k9IgD0UOinpFoIZMT3eTaxyQe/AOGkNGjgKSxEFPChxv/CF8cHKkXboDsg1/kyCZ+CYdNOMEMNhgIiSq5IJYEch2blM06wCSMv/2DHojQQQtbyEAFrk4i6EgFOhIzuSg2cy+M/Mj4aBfFKHakaZARHIlQqRDXAUIVYqshBwkzz4HoUzOBhAguGhqlFQ6GBzZwwh9scFGFzHIhBWwit7jpRIYwUghSqOLOsv+ZykypIp+iGyRjDFfPwkzxkhyh40ASChFibsSOeJxIM1wDUY/wsjBnY8XEJBrUiTTgZn/4hy0GAgboQQSb1RInR/7JkyRAwqQQxWlS9fLBeypUIQv94T8e6sabujSofvyqWyeCDTMs5KmK+MfNJpKEJHxzQXpj0jf/KpG/JWETK3BCbRbCgyr2lUnCjEgq9Amy/b31IyBLxT1byZD92SEadtjhLlenRono8h+nIO0pYIgLOADTU3Do7D84+5hm6PMHlYVEaXW6EFZIQxdIVUhbT6cQYIKMjkOtVlOdOhBqSpUheTXDNJ2315X9Q5zPjMw39fA/5v6jujbohXed0KD/f1SonrnaCAwF4sOFSANk+jwFUB8SPq9ChBXFnWx5I0LM8K01AqnA7D98yIr4RaO3HoHDNOCA1oHg4qHp3ZZE1/ANxuTzv58t7Wr19w/XwoFrJuTjb1VoB2B6y6YPiUaB+GhC1yrkqf9QhBkqRFWFZDUcC/EuO1iiVyluoroeialE9GqbDCnEqoddSDIYYYbwkmgF/v0IK3C7P8mmwoep+MEpSruQyn52IM5oMkMabGLcTpYjMKyfY1+jkPRyjcAe0dojFDyQN0/El1368EYGrGKGYPkfj7gylqPRYIaw2c6CJrCJMzyQPaPHj9ioJnIVYoZwwNGuDCFRN1bACO8yYeIfveC0QjLdC3Z0I8cTWUeMNyIMegziH4M4zUCemQknJOMf+fj0JDvjigqdZhDOqK9HGswKQKdhf6MFGSsCzQ2j6rYjaw42Lg79VRJG4L4S6eH5Es0DkJW2wfGLcJ45EhAAIfkEBQoA/wAsAAAAAPQBGQFACP8A/wkcSLCgwYMIEypcqBAOw4cQI0qcSLGixYsYM2rcyLGjx48gQ4ocSbKkyZMoU6pcybKly5cwY8qUSYvGwXLKBlYTCADApGqTelYDYMFCjzu5eHHhNGfOzKcMufzjwgCq1atYs2pVmEDghEMGJxncabKcF4HlBAIRWKJk27Zb48qdS7euRxls/oUi0sPLg2UI0y4UAIDiWYGHM3pRNgIsNIGLOsK1S7my5csxVQ3syaLVFIiHy5Wz8PmmF6BDfRY8hpa1QcAGXWfsgYAT5tu4c58ZGSk3RRCxehDMuZCFIUN8RjxYvjZkOUzVMD0QqOwB8Z3P02ovuPgYpn+FC77/wOH7IILy6FPG+WYyQPqFLQou+DciLfGHM/4FmjL9X87/DD0gGEb9/VNggRZZQMgva7zn4IMQQmWCR5A0oIQx/5RW2kJptYXTTQOl9ZmI/5A4xQ7BGNJJcqIFVhCC+VE33RQjZDjgfTkNONAbvtjRQIQc+QCkZXEMKVN8fhDxAhax1JjDFCUskdCGByaUCw7iVLEDQVWggUYwVAwETBX/3FKjYA/Q+E8wwWy5pSECVQGMIk38U0UwaBgyAxrAFDLEP8DUV1Bz/pU4kArPBKIECv+gEEggwTwjkB3WGGnppZhqdMZkuUww1RMG5TCQqP/EkkuGC9HIx4ZoBVNFE7fc/9JHFSOMACYakhhAZwgFxSroFMEQhAYVkvxTLEF99DHGLcVWMQQZtgwkCRlh2mpJCil8OUVparCw7Qi5BCvpP8/E8eNAeJCa6bqYfccuSVxI1cIMNf4zw6n0DeGOQHWOoEYr/xgywmdqCKRFwVPEIs4thSTESEHvIAQOOf/0Qc4tAt0SQh8hdNNHnVAMNA9BIhDkD7/FDiGJJENQQYUhbQYiUCdh0jdFOVMEUmuNt/DwI3vvBi10e/8IsNUEVXGRnBW1UmGJAUEY8HQQwBzUsJgpSB0LQWpMUYWsBfEgkx3/ZPKPDS0HIVDNKWTxjwGG5BzIGGvcI1AD9gxk99B89/+d6SwM8ELvCDM8bYABbyc+ETJl/jPGGCFsEUIMuuhCOS6sWHXF22HK0zJBVQs8gqJw3NNAPf888g/qe/vt+usYAVGEQFvONIvS9AZz7eGIGzAE4gipHfxKuKBERa1TGBOIj/U00CDs0Eef26mzCD7DDJ3wEmYnBmTN+z+/H/4noGJeqjbMU6gwAjm6NOD8uQOVUYb0HcH/DyT0m9SFKP/IkmkHRBAHH65Xghq1AltZG0IKxqcQYEhCHDYgwD8wkAkkVKAgegDJGI6lMioA44PAMEDVqtbA8jEEDf6qFfvc5757ZI4gBMvfbQTwBYK4R4bv0YYAZ1CC6/GBFwtMQQb/EIiQ8YljCFs4xTvO0ZIMEmQFaCPhQIC3kSAEY2cLYqEq7lCASgiECQJRwT8A8Y812I8g55HLHgQCKhwy5AL/gCNK1uhGhsyCE8wQXCtmUAbsCfGPQ8xARCIQA5icTCUGQOHOqhCIZ1yAEnuoxCPhiIdU/OOMdcykJjnCBTbwohVlGGArDpiBLGSABIUYw0KcgZkXFpGKEOGFnmagBh62gBKUuEAsUNA+9zVDggPYpFVkI8zc8KEDU5kFB7RBiT22gg/B6MQ+QPEPVhaTIFlDw/UINwI+5IIAfpgF0iZAzgn4AQtmbIAuBGABLgxjHO1oxwHmKU8N8I8S18yNbSSC/6+VSOUftasMwBQyi300kw+jbAUl+EGHP1jTJTGIQR8UoQhlIUSV3cCKIAWy0RTsA1tB0ObgulaOrn1LDbWagRVmwIJYzMClfPhHTIPhzW8agxwo+AU6dLGGCIijIGzYJ0P6KRAftEMgGphLeD4iRq0IpyBttFRhemMSce6DF7EowSgpkYJCkCAZMInWP0LAq4F8Yqyb6IYtPnHWf7TVrZ9QxD/AsBJ5bCQFikuIIPdhiU6waQbODGX8SvVSPrRgFn74xy4u8QtfyMwCBGEBE9oi1Hxadi5fSApCW2GJDHguD3nog0QiwJFDRuwf3+CVIj7hhBV8Q3XYEEjx6voSu/8K5GoDcZs8MrCNDFzVEq1Aw5pmEAzAxkggwRrgP7LHi33sYxWhyEM88mk0giz1sgNJDEsA8IYd5IISyDFABo6QhUKsIg//2IRWVDfbk9jWKmIQw0Lc5rZ/NOwI/9hGFrYhj97ydxXayMAhVjEMDWigHQY2sERMsYFLVSUmT8hFVLH7kF0I4A13aAEfDJEC/ZKXH1l4WB8WgAQKd0S+/FjFKq7AyDcEYgeEWEptGMAJDnCCCx/YgQV2sIM3gOANb7BALC6Qi0jGh38IeYOJtxLMgYzjXaBiADTYoA1trMK54gAGFQzQ3CzIw8tZaEMbxHAE/B4Bt69rg0vwe5A2QAD/GXnUMjAsIQ5xcCEDV1gFP3ghjqQcQhyJsERzW7APQnPBD4HuRFLo0IUlOzojtKBIYv1gUEp0ohOtMAQl9pEF8nq6vPXFIQlIQAcSCIQEEPhHqlP9ElOb+h/IWAUE3owMMfDDrp2gxHd5sQpqNrrRKXnDLiwiM4G84NHvAQQZ/1HDHcSCC5bggjZu7d99MOMf/EiximftZmQg4whk/keZxW2QUP8jHxFRJUzGUOKKsPoioKADFOgAChLk4dUEoSZKkKHA5vLCGDs4ihty4YEEdIUyjMrUJf6BB4E8lSDVVQgRbmOMKETBAsfmCB5u+I8P/EMO2+CEikWwCgWcNxSr/9iGE4bAhSw1wRXCiEAznNGMCjjD5v+Qwj8qgAQkqNcJUBmEQbYRkTaAAhSrEAcO5pCHWFdE3xSJdx7QPbJ550HF20DGNgqxDS4MAUsEeAYBxk4AORBBDhKUoNEabrSF/wME/8i4RHyB7I+43Y29oapGMPAPPUjhgv9oxs5XIHSRwGIgNahBEuihBycOpBnnSEINFuIKJQQCB6tgXEEYp/mCpBoZSK+CL3aBh8Uq9gyBIMcz6rwNHHB9G9vIA9P/Qe9/UHMV/0gAHdBLh3j0/h/JoMM/8kCH3vc+D4zgxDYIQI5hB8A93mgEVQlBAZRw/FKaoEgcikQ2IFWKII0wSP8tbrj9ZT+IAtRIgjAqAHjB08MV/xDGQwkCeD0I4x+T/0cSAK8QJhrE/wYheP8AgNV0QfCnBAYRBliAATdAEKEgEK8wEIywCvg2EL22CulABzeAAkqgA4tiE76gA/+ABQOBBST4DzaxEGZwEAg4ELVQdwohBCahCyuRfSRBRuZ3Gyn4DyJYJAkhgmfTWsKwDltBgOy3AiuQQeFgEIIwEHx3ESdQEFEYhYgQIZEmEMXwD9kgTD/ShRgBB2mQBj6IFYCADpeiCuiwAq6wApmQBHbBfwqxApAggjIIhGVjEDYYEVX4EmY4EWR0DZoxEdmgCoO4hSLRh5oRiAoRiKpgSTD/yDdwMA3/IIn/gA1gQFcFwYYGkX8FcX9aMYRP5AQiYAbUsHMEoXOPSBDtBhHcQBCOmBWnNRCqcxnRUDyPQIkgEQ2X0SDOYANyVRArGBE28DCk0Au9QBC9wAi9wA7soAgr4IkeQXiuAH+LRxBuOBDodm7/0A9m4ArUQA39sAKLlwQrYAYldgpulAauSIMkIQ3sqBDR4EoaIQWk9R7SkIr4mI/6uI8GMXHPczcJkQZ6hxDdV0x5KBBJw48l8Y8KORKJEBw7MCBkERJAQR2QVS8rwQKR1ZAcaVlzAF2HoAKTIBiwwR3/IBYCgZIDoZJX8YAd+ZKP9kIDKRC5sAPVoF3//1CSEZEj/nEMOqIQiYGTGLETABAIfpAX/1BZElECcDE/MPmUAxF+L/gP4XcpZlgYMlMj93EQy1Ad/6AGNJULM2AW1EGR3CUAFmZhArCW1UV37uELzxcAcCkAchkAdPl8AhEAKHADnOAB/0AA7QWVlxVxA8GQJiaJIOAGOzkdapALhmAMOGEdOokZO/Bngll3mFQSY+ggyHRJqfAMTVUoEEEvOGMdheKVD5ETO4EJyqACESkgFDEiF0EWWMkgl3mbuDEhGVEJYCEQJIgBEbAAz4CREZEWOSAogTEChhAL24FcwfAZI5Bp/yBcwBAs/GEQhvBiqGIvB9FSOaOcWTMw0/+xlSGykpjwBr9wLnZzLu6DWv+gkbgZn7exAG3BBBqWQmqgAgVTMP+QA/yJKnwQmg/xGTlRICPwNaJVBd8CJwRBLAMBBlcgDvWSJjViCC/jJXGCBkPwJxjToFTgLJLAK8UCJ11TIixgCbHwGY5QEDnAAmKhZPrxDxQzKfL5OmYhlJc1C//gKbcjOALxnwOBIQMxA9tSEF3TTVUTDF0TCBUoECOTD9mIENigCzogpMFyLAJRVn/wD2SgCH8gCX+gCBD6D5tTECEwBn8gDh7EW1r2mFPAn4YQUinyMuJAMc/TIIZZo3qqEDOpFRNwaHzAB1SAIbmgZQchWqFDQn61HwL/UaQ08gy/UBDVBxG6gAu4wAM8sAnuoCwLwAOVwwMF+RDwl6UhgDGKwA5po0iWECZRMxAfOhBhUEgCkad7Wqt24UVcwAFckAtLQEtgAjWw9BBytTJ/0gR/wHVDUAVkUitkkhUsUzPCIyYvc6Q0AAfuI4mqgzr/oIi22q10wQX70Aq1YgyUcDhZ8zbjE6wRITYDkTlkUzyhChMZEATbIAYMhBDHMwIqYAy/YK0/0jqZ6a216h4lOTszMQCzMC/0YghA9KHAkDXnCjuWgEI00gMnwEIHMRkCa2IOsC6IdT0zoCL28jQJ1D3gMxB4JRApW0ICEa23RRLsIBKWEAS1ogY9/xAFqcBCXcitqfgjs+gSeuceObixGLENh0BAPgRE2KJAf3KvA2FEkoAESiQQNXcS60APA5FBTuQKOBBCIUGz/nKzPpNOWyRHBAFZRBsRhXFdWKGYceRos6ANu2pc+XEt2DJETPsPK0sQ44MBzaAH6icTN0AGh0MScENLhJMLqtAArOAJBQBJkpS2LuFFkjsBHMAM+7AHe9RHurMPQ5ABoLuh9LOyBkAFSkovnNUCewBJucQCXwAO51KPB+FxAnsMs2Owl8m2CyEkGHFHuopQxtUJXUUCNhAh+DMSKRBSO1MCfFAJUUALddMACyAHDDBO5mROYeAQDaAKeJBxTyYQB/8wEELCAJVwB5KbG/DgNzRmUEzwTFslD3lQVgkhuyUhq3WBV38iRCprAH81UrXCB0/QArxADnGgC2kACOzEBbLgAAbmAxpwAA+sAV0wAInwBDqwBs2DsXhaEPSbKbprJERFH/+Atv8QBTKETwJBRwcxCwkbqAgVDLwgD3SAiSpBwwLxCaTwVgahw2dlBC6xUQ8BxCqrOMAQBFQQUtq0R1dUXAPExMYlSnz0D5PBB9nDBY8RVAZhEySsEEf1D0aVVH5pqxPGEgFFEghyEuKUCyzgB88ETdK0dcIXE4eEDX/wViGADbEIWwIxfyhhbiCxsoJUXxlQCLxVyEMEN84EWP//sEdQHFOBikv/oAKS/ASrO0ktMAfh62g4er4CsQsAYAyWkAumYgn6VQhHkA9kIBDzMR8wEVvChF8N01uFkAWm1Fu7tQ+gW0q6bErMkAch08USYRt54QKw88EbYbau45IlgQdv0AOJQMVd1WlZ8Am9kMrvcjX1JV8wwWYDMWbehgz88G38AGvj1nmdp2ddZwDK42wRdgGV0AFzIAoGhmAaMA4aUDJ6OsZ9gwr/wM8dkUY88Z684JiWgMuz7Gnj1gvFsor/wMokwa65oWYeoWbdBs6Zp2LpgHScwAkIwABLwQWEsAM/9mMWAGRCdgFwRAlckA4CwT+iwD8dW2z/AKOc/3xNG60NLCcO2wANGWAJVeDCvJBf9EVeBqFeHxEDfBwX7yYQpFAQTfoPT50RjMNqq6ZqBCEPKWAJwJALlkAJXf3VuIRLuaZQipYL4sAJXeAADtAF+FzTJ3F9WlEk0lcqfsALh1AJuXAIsWAMh8AMnKANzJBHvCBog00J4tBhZVZmnSYPs9wwV8PNqmgZMlgSoJAP1DRqJPAwpzYQ+BbVIoFv/NbVSsEMfsAJKKcNyjwQW3wVcPd2bg0R5hvbHfEG52kM2wAKeQABqIbZut3br8Y4YvYPEn1fsZYHV1AIhYAMyG1fmyO/vqFeW4DPncfZF4FeAlF8ITMyteduBIF7A/+BXleXclUAAiBQemhZesP2D3yd2geR3nT3lG6XcBjxASdoF0I6Ep7wD5Oaxf/gCzTg33EHd4RAAOtnTfNXATVAeCaRf4c3EA1uEA8+ECWDZgNxBBJdEG3AOKCAA7vQ4cN2A1dwdaqGaghBTdYdESY+fAKB28Nnby5OAuelYghADlS1G/qddgVheoolEA0nED/1aDRYJJsJJDhYlQURALUglVlh5BbBKBTgCuxXc1Jwc4vXhiuQ4OA4qhMBCzWAtYEngAL4Awkh5lQrEBWwDoknEOYwqen9lzgACnNAAtPdzcJ9EHRQCIGwCyiAegPxAmeAAimoBBiwgAWBAYyycO//bRClWIr/IA6eAAI23igWMZUHIXcSQelGUgfpMaMyKhA7mEmIsIe+cHcCUQc34AqZYH8rQA01wH6mCBEEOBEzN4CzfhAPpXORd+UrsN8CQQ5N2IQCIUEP4QvF4Au1cOwOPdkuKJg8SxcOQRC4SBeAWIYDYYZ9yBF7qBKhLhCoeBBTuAVmII70kATXWBfCkAnh4IaAtwDZjgRCgATAblmGKBJX6CABexG6eBBkdI/ximxOELNgsITl/hBEqBXX6IYHqXPttorQSBepMIZDnhCqEAfXXhEVDxI8+4oJAfEP0ewVcQr+gI7/QOaXcQovxArRIPIfEe2X0QDhELP/sKUC/+EErpBRC1EDtmAD4bACm5AE6zCEDS8QQa8R9yd5P58QNZAJNnCMTc0IycAI/bCEmWAG4YAEAlirEX8RlqTxB/F3D/Lslv7aYj/2ZF/2Zn/2aJ/2UAk0BEGcBSFGLxAIvvAL4KALDiEOTiEQB5f3hBk9/6T2gF/BxqACq60Q3zGRY+EFXjCSypA+T6AUL9D3KyElGpsVgAP4aI/4xKQRiD8Q1/Ge3An6JDEZZVD5mH/6JGFy0IBV5XCT/7DJB8GSKTEClIv6to8boRCSkzAdP3kQm4+SqNESuhsZkfEPxHz7yA8TOZADTMABftADx3DGFJEW1cAasH8ShVENbmAbLv9w/BYBA/8wPzJQlslf/gpBmEuQCypQDtPRH+QpEZ1vxvB/CJyAlOaPbJHmDUHT4yoAELGAlCP4r9yyfwkVLvw3ZQQfFtUYTqRYjuLFf14SHpyoDOEyZQqVaVw46Z9JhT24sFm0sAFGmDFlzqRZ0+ZNnDl17uTZ0+fPmI0UChUK1OjRiQCmNFxKUwWfhLF2HHwAEum/Y5gk/sP0D8BXAWF3hQ37L0CAYgHMFmuU7R+4OOji/EsDB84COQpTXeXb1+9fwIEFK2TVN9JgxDV72Cw3hY8hQyMOhgzJF+GDfwgrJsR88UHlhMcWCvhnDAeBxKkZINiW2vXrhahgz6ZNO4r/Qos0R+TiI7lzQs21eUYhEGGNcKQc/ilH3tx535eIDyc8/txomIRwlCy2+FvmjFiNy4EGzTP3zKaNfQJI+OxEdevx5c+nz/MLQ7X/4Nc2cTVVAxqMSagpp2aQbCny/ikPpt9GMCSWpc5bcECGjJmBIe9m0mgS9t6oBY76bmLuKBFCNPFEFC+Cp7+rWOGBnMWmWIrA7ySDaYruZhxwBhwbczCYf3I50CCFlhqhoYXKEZAhh3CcIpjIzpvovNze2EWXBu5JcUsuUcyPtH+m65I+P4hAQYgoVEBSTTVoZAi03zIcMJgqgGxqBDSCCSaQYNCoIiFghhCSImM6McRKABoD/9KQf6hI4Z9AjmR0hGBSMOCfYGzsaKJqQPBljeNAXaOBUb8Z81RUYfuyqFRfYyIhLv5pIZFEDqmED4hYUGEENdp8Aio3E5oQpliquOWWKgKxCMgq/EyoCmASorOKI5Es7R9D8lwKyH+q+LMQhVJolgo0HJXkFluACcZNR9pcKEIJvJroGRRA/GeXVvPVd199S5DhnxIqaSGWav/JQaGDGWqlJi3+AcJhhTCL5Z8++kB2hClmYJRcaI9g6NhqywnkwoW8peIfSZqYaAiFDDiXYpVPbojSFCwxJth/RoBwIh4UioZfoIOuyS2JJkFJaMQKSGiCCWbhJZZd/1FzIUv+Qf8N5yJxjOWCxYhsdAhJbLHlnyb0rALsc2/5OKFAerBohE4ScpSiEPro5h8eYmgC7EsT6uOfbvoQBxhDqKAigxSoMIRHNf5pfFA+ZO5WB6Qrt1ymkEi6HLFYGfhnlkRYYCGXXFpRQQ0+yHiLbYV2bpxCGXP5swlJWM7jH48VQgZcjHD5B5t/nsF0CDJu+VuhPkJogpGFmGckj9spckLlQIcwIiFtrV0omFwCAcSOURsQf7/Nyzf/fL+4mCAXh2bIRdogEgL3l38oEKc0SrDHeCEtZOTjmVs0gQxXwEFOeFAY5HUjBIEbwwJ40DOcKOEfLEtIFqgQhMjsoFGSaxRkDKH/J2NU4Rl7CVV+0HdCFCbGhCaaRawOYQlepCAF+8jANjIgjxsOARkxCUIuIrOQNo2AEOSg30TskBBd/MN3MMGFHZq4RIZAMCGoUcgfFmIHXfgDCRH4hzMUQYYhGA4NhojfP4LQt4SkQBxVAMeoJmKqFMZRjoIRys+ss4d/TMBzvGABrxxkgDPGLwjAiBbKGEI7uSWEZbUDBrUwpoYRVIEcz4lBGv4Rjn/8IYxB4KQZUyAPYJzMEIGYQiBoEL5QLaQYRZhjK11pvll8zg+9OVInLAFIhRRSJiy7HspUtpAmVEES3XrGGHiAiyTS5oiKDOOlWPYohSgOYyMYAxzEVw+G/zSAFq/kZjeFxgUuCGkElDJAOS+FxkvpMiZHwIBCwPHAGOwFby5KIhR1ksye1M5S/8hAy3LZKIypgBxtjI43DQoU8h30NbPYBx8MNANLWKqc+0SjTo5YGHwaBYFHKeNEohWEcarBGKck1US2qVCUpnQhD/sHK5szixbMoASUiqgBLvgPc3qTCpbozRR6EIj/1CM62FRICVR6VIOy0qXIucDneDEDqHYihn2KoU3RUNFXRmYKamCBErJUUqKqIiFGRWpZzZo0p0J1BrZc2C0ttc9wwaSjmzNEr9TgBh2ErwFETcUdzrqTlxT0r0ZxgEJEgb4JbMMPsSgBVI80g4kawP9SFLxJIdWpOtWZwZA/OQVG4qdLdf4zWqFdyGhB6kdjLEB8q50IVAb72tk4oAul+Edhz9cBNxzCoY79Bx8iOgQZGoCyGAGGONwRAVycwnfvEEw/bDAIV4TjBq6YrhnIII6q0YS0nkUDr9QQCxR8Y6/i4wEhKGIBhWgJtvGZyz8AYZR/rVcwTf0HMw4RC976NgXAlSFwYfIocQiCB531hx4EkwSM1OAGQ4gWVn0Sre46JBZK0KsqnqE0hbxqagohqnzj4w0Pb2kW2uBFLmaw239EtL/73e8/oOlihgxhCz/4wWtqgGBhKGQQOBhmXx51WjWUwBgxEF9fC1CJptK3ayH/lg97fILHv0CZyZ/7BxcoMYMynPgfUgUu4oD7zLgy8x9koAZyIjCKf/DuL4DsREhj8YxfpIEclUByJaSMhylXjr55DgwDmNHQVswg0K2wxD5SgLgMDKGfR23zCKxQgickYg90psQFKvEPFuABHILlc77e12m/JOIfDOACJxLh0EEbYr+JHsIRmBcDinCxxnIcQt8M0IpxQpUSu75Ar2GwC2mslosKacE/BvAPP5j3Jgy4NKhtslRny4cDs+DELK7sUFxVjx+McMc/hr0QLjrD26jyB0MeRdnhUoRlww1Cd8dZgla0gBLgxZL4pEAEpk3AD8g2KU240OxoY0Spogk4/03s2BeyErvKHJh2K1qBqxmgwRLbWMUvv23WRyUuU+PswW7O0Ea8MECPE1CfvsMQDfGh4xIg+IcPNNCOdvzjADJPyGELntIuLOQV5itBLIiwEGaUGOIO5wUJ/rGAmVycPs2YDSD1NIIZQLIViWgBTGGq7zqETxfeAAEXRCEKDfjgAPg4gAbK7gAru+GUcGSIlmbdrTiCick5v8kbKrcPhwsaKrzIAxgoIoVxJ0TpRoF1QiCBt38UPlUGQMMMNu7dEThiBCoIxA4CoYLRZYAZ2oDGHOaQhzmkIx1zGAIvKPEMaYxKr/eITo03MEcnt2oDppDJQyhSBJZPOZZsCKfj+f/Qik7sAwLMe00fxPYHRSTECEb4RPMvcj1SCGfRGMlCPw/tYktQoRUbh+RWHQJJqKvVoY1trFr/QbCJxaJYhKiCOF7vAoWw4eZ9ef1MXDsR9Jb10/+Q8kLAOQuG6gRccThHQYY8sAHhIIVPgIkFJIVeiL4tGS5oEiQzmojgsgQMCjSoCgbxA49/WJgsg6onoIR9SAgOuB+YuLRmk7+E8IFWipf5GIFXWYgnsBwvOI+jEYz14QVeKIFg+L1CG4I8YIe7GYPaeIR18Lt/+IQ/AJ5/eARs6IZwcIKE+AQwGANsYK7BWDR5uArJwoguTKMg6IQZsJBAg4qFSYjxYwE+oAT/SyAYhuADS/sHJPuHOdCA+eOXfdOKzQGBJ+iAX3mCVuCFG0KGZGgCI0Q6mnCGCFDEnniEhPgGI1xAI1CEbngESJwILXwNNQsMcAlDitgHXsAgDgQSh/qHE9MyhWiFXTM9SqCzCyg2KBAFKFgIPMzDU9mKyymCL9iBROANVuQFHCqEPLgCJGAIR7yIwdMJbFgi5nIGZ4iBb3iEd3DCVgrDTvyH1uAnG/qHfTA0A3BDQwg0DlwYbjGEqjm0fRgCfgCFf3i5hBiGmeAEXGwlgoONXXiDHuAFXAm+LNiGLLiC6KEPKDSrLDhIhMQhhMyAQqghh9yGI0gHWdAAs7vFmzAF/xegvVaSO8DAsJzBRQB4g1zgKUvIgIMshCygAzDYhDnqxCwQA6SASZ7YIWQQA5pUiAVMCJnMnW5MCIrjh20osSfIhUSYA7B7OYocB4ukCXqsHAQYNZngyMC4gImRo1BQiKtEin1biF0YgRZ4jBQ4yUI4gitIhn9IxDjKnX/YIX44CrW8CQggAVDYhoYEyG0Ygm24gjlYBQVYhQRYhVXYBnEwhkB4gx3YARDYAQuwgK3JhQIgynQYhq/Dw3F4x3/wBF2sR5mowTzUt3+wO18QgB0YyVgIy4M8giw4AtVUCJbUzJiAyVUABQhABggABX7YB/XzA07YBk5ggN4UuQ84zP83AAHDHE7GHMoLyIUJmAhRoK2EqAYNkq/2AgRWcU2biBVF+ocPIIAYsgRD6IRDA0h5kAd+UM0sSIgrSKk2iIn1NAqP2aGEaIM2mE0Gy4AM4Ad+WIV/oAP9XAVtGIIqeAMBHVC70yCoqEE2iIdXUNBX6EsF2DmFwJcQsyTrtIlj0wY6+DzA5AdkUE2I5AcIyE8uuKAuzMYKhYncac/1nE8IgIAsqDXTs4ROIB1L2DXS6QRKwNFWKJ0PLJ3SmVGKk4V/SIATLdKJeMpj88V9KJ1WQIOFoQST9BiURM23VMJjVCgISI0snQgI/IcWhYAjYAZLsYQatYQb7QQ03YMcpQT/XpiDf6A7E0GBF1CIOTXShLC7+DgpASgCaGsIu/MDcVjOz9EGThDFGM2FndoHeQDI00TI3DlPhmjNE0nGvyABOjC6uNzS5tjS+ZzP8kycGeUFbQiFBFCABEgACI1TO92S90qIfSRTHuSF0uPBFOAFcYihWN0GMWgDfmgDMRCDIwBWj5FS3EkIUByTYzTCxKADOsiHfyABEhhIdzQ611gFZEAGBsuFGeICN+hWTkiA24GHFMm9FLqNv3qvVv2H+wgEXvBPa21RElgFEsjUeZ3XL0UGX13P1VSIQujCI4CA9jwCE3UNTOILIdjPq2DWfGBWUMgDanVHndBUL53YibjW/xoCUAHFAwHtgTuoSoaAhxIZjX/whX8QABRY1RPqGk/4hzuo0/X4gjcgjV24gVVIh4aVV3nN1C9Nz3+4gvyMyyvwgBsAnEzIhBVYgT+4ATIgAycgRka4G31h1tuJ1x1aT/jECXeE2IkwOq1FWDpoWIzYUtqk2H8ABVCwWRFAAC4QhzWKAgHwhQAYi5LNiUsY2SJ927q9BBqYP9SggG5JFhrAF1/YhUsY3DN4gTMgBApAgnNohsZVCGeogIRYhxr4hxpYAcCo3ISAhZzYRoy42vVchTyogl3whWcYAlDQzyuQ2ISg1oXQ2oHEiTyAWOa51CtYo0DYhbM4i0hIC3LYTv+r+Yf7oaJ7wbO6XQhzRVmfCISZULajwgKK2FuFqIWEOIOTPYMb2AJncNx/ADzJ1YMaGIRBSAhXAAzOhYUaQN9/oAfN1VyMoAYqrNiEAN2E0NR4bYJdoAEUGItdCARxoLjPg9a4bF1G2NLbid2EMNuLgNjZnV1QIAFGiNfaXIXbfQa2+IdiSAjodV7UMC+1WCGcCE3lRRXqfQ6iaIR0xYmT/Yc6EIcVOIcKgMZ/EIbwTYjxHV9q6IefWAF6oIcKqIBmYDpneDuKgGH2ZYjxpQAJ8gUdKCDbXMt/aMux1Z2FmM3UFYfSHVxfUALmlaAzYAglqAJCIIAPoADFJYQwoAH/uA3NXUABAmgNDwiFKxCBUAiF+K0DSFlhljuMWmgEocjghHDemvhiZ0ui9kqoyqFOQGaIbbqGFA4aCnCFCtCDH04IcZvkClgBVxiEdVCIcxAGBEsIzGUI9A1lhjiHhGC6iSDihdjef2gGyY1ceviHfvBbu2WIP0lP6FldjHDdVfi8IQgDFAgEFCDke7nlf2gnhpBenVjhnaiFEsbgsxIEfgkDapavk1KI410IalgBYahkPcgEV6gBPUBlmYjlLroIIL5kn0BlKRCGo12BLZgIPJ6ihRhahhjj9qMASSAASRiiQBgDFFCCgR7ovaVeyqln6E2Ia6YJfP4rWviFbB5h/8uJ5om4ATPAAWrIhEqWXHO+Cclt5ZloBnHDiJBWCMldgXAu35yYZ4Yoon+A5oTQAWZeCMqxjhNwC56YaOsQq1OpjmXSF58+Cpj+hxMo6r44AYZABIzQgbpdATNYgUxIkU6ugCRwhUwwMIVAhIPVBJvg6ZpQastxi23S6bMqqMDKCRCxJHlaCKb+h6EWjLh+L3RQiPbyiW36BbFGDp8WAjMYBFOe4YXIsU6ejwrohhUIaQTThMPDiHlWZpjIhrhOiLd+jbm47H+wBoygAbFSheq8CclOiGwwa584AVUg7X/IBnRQhbqGidZGkbTmCWnACERIhbamjYxCmi1wAieA2v+7mer46OQcowkapgClvul9SYW7vmuMEKtU4IZ/uIaccIu6Hu3XPorXBoTJxojVTojbpuhTObhogIPx/ocQ+Ifk+wczCIcbs4nhlo/3dgVXWAEdkALAaxWkDpEr/Yf9hgnphmu4/m+e4KIi+m6daGyhQXCM2Asp2hw7aoBucIL0VggnKNiLuBsESwJQFux/OGmFCGy/yLH3Zs1/WIcVcAKzTAZ2wGpqcAXAQ7r77l6K5obnPgoISqLrxgnfOYVMPIWD2xJ7+gdp6Ky++HHYvgdsUIQJXwgLjwkzMMuE6IVkYAQnWIFu2ARhWAdhAOUcY8nC3uEW92YOXwgbMMteWIj/ZKCGHKYG9l2Bblbl+ghy4bDtvqDQmpht8M5zPd9zPu9zP/9zQA90QR90Qi90Qz90RE90RV/0PU9X9sgP+ICDJk8IIi2r5SQ5KmN0TY+JvLKXiZCAHqA8xZwCFdgBGVGB/CNmFKCB/9VPhriChVYp7KyyTSd0BagJDFsSC4hOhtCc0PgHichMr5gEZVAGFVABN0iEUlsFTkheszq2Whf0UsUIDHsCXRF2o9AIbS+HXYmC+0gMPFuIJZCaaC/3EBmWv9D2k1CGgjF3d0cfN/2HW/8HBDgEUVuI4AgMzcGM4MiNEmABxCiBcX93gh+Mef+HUBiAJ5gCX1eIewQOrMgI/2BHjISRCfgreIyvjzmYd204hCgoh4bHiEkQjZAXDIswdorgBA/IeJanj1sPhY5XgUmwiHyfCJOYeYbIQcTYiingzJb/eevQggvQSGg4BAuYBDmZCYn4il+v+SmReIkoeZzwAhXw+Z8A+ISDQaDfeprggFAQBxV4AMyQ+pn4Ci/QdqdnCIsoh0mQCCnpiXJQiddryn9YeZuQ3oTjer23v6cBgIZPe5lAiGrwgmMge9yAeomHibeXidFkwYTQyJswKsnfe8q/CIDfgbP/CLhv+xu8CJTITJ2PieAAfIVgD2MYAm1oiZbAibyvfNdPCDWw9nLAjKSnCC9o+824/YQwGv/NuEHCv/mHvwmE0AjSZ4gd0M1/4AS6f33mrzuC6QyQX/zM4AyDGKcNm4hlmASNcDIBYI9qaPvP34yFCHa1P/yZII1D4ITVb372pwkAgJrzeICQz3cJ44Ol6PyJEI2ad/uSAIh/AgcSFAjg4KRjkwD8AzDp3zGImCI+FPjwIcOCHxAU7OjxI8iQIkeSLGnyJMqUKleybOny5clGMGfSRPmmR49/ykYu+/cgFh9DsUZ4ebDMaM2CBwEICECw2L8AkYo1AgQom1VA6OLE+YdOKyCuXLMRYoCA079TSdeybev2Ldy4cj3KnGtXZN0eI3b8K6dz5BQ+QQOVO9qTrd9/Xsr/Lfayc+CkapGPVTPY8LIAAR7TNCLE8S7o0KJHk1Z5JqnMuqVFW1A5QqCxcoWNPnCbuK8XgUj7CsztkfEDL5g84jmENtXq5MqXkwwFjTn06Gt3/Xt9O2TtKTMMzZhSVHTiZddN+o04cIcfAtJdTljvPiWqUO87qppvv2MgFgPH/67eyhBhR/nUk2/3eQSAGxRAYqBJXBDEAYMROvcPKgLJ5x5yETLXQUe/GONaKyPIVqBPJZEInQXPRKDhSFxACOE/n7E4nwLrNWBXJDOaJhAcKMQyxUmy8fGjbH/V9hh2iflWmG4ChnbQDs+coCOVVVrZVo5dXTkSK2eIGGQ5M6hQ/84DSNZWG0k9jSiQX2iahKRu/wChElP/BELDjVsSxICeffpJkFR/gtTACZ6MWSJJ5QAxgxrKlGnkXympMIN1A8HZ3xSBGMMXSjs9gGZFb9CwhkjSRMjAIjX9ICirra5kAk0cQtLAAjkJNGeiU8SiRpEguXlkiZ/6VM4OQRkyBX+83XbdDMF89MBtuMq5H6IG1bJGnh/B4apJw3D7LbhwYfDPGuS8BqRAWoxUjjIlHJpsbW1G+s8UUyAZyHbBADgevwTt4CxBfjn6zwwzFCmttOj2ttAuaZAKkqnhSjwxxQXB2hJU/3DzTxy4pEKOCtXeGpJfJeTgF5Bu7gTkCDmwKf/QDgUDOcUIrQSDRjBUfBkwvUO56RFhI4yA7AjBGNDJFA8gzNtOcB6DAjrZCiR1xVXrqZnVSfnxz9Zb/0OADidsWpDCHiU8b0c0V/HavNzRe7NAVQADDNsj12sIH4FkVF0wzqLxDxUCCabGFMF0koE4wXBaNr28DXQMCOiQ+vA/DVhOddaZRyiAapqzx7XXW6Og6WNAqtHRzwI17es/xhizdpx9o1E03Ib8I0kVtyTduED4ChWIALsUPpDckvwTzGt8CE2FOMBUQQXjBa3+zySB+IKOLqnEsdUvvyyQoefhv4e1+CntklMJBXHBCxdeE/JBLizkoIYagjni0aVoF/T/gBpVkFFILgqChgF2pAnBqEIggNU4NBhiL28omkCoQIUhNOEfckMDFQaIBgMU4h9kqE70PjIJob0BE28AwBt2EYhA/AM5lCsfDKHTuRh+ZA3U+Ucl/hGLEvCBBSNQww9VoAYVTIFw9FIDE/iQOpKkbCBqMEYT3HEL5NkpKH/7hyHQIDdkgGEIuNsByh6gnX8w8HhYtOAtJNFBgZBhCFWoghYneIs+CARg/1BXYIb2M8aMQAWV+Uc1psCpX/CIhoY85H1QAIN/lOAJiWBByOYnkNMNxHQCaQUlR3K/mVVSV8/oQx9u8Yy9OMt2gZNbB2/xjxDcogpl05cpzwhHA0ji/w+3+MNA3CgQYEiiCXSs4BUH0gleDO1+BbEOX1jYkW0hspnOXA4KBFIGgbSgBe4aiRqeUBIg9FEZxlQXvaogECki718W1CIwhuDBf9yCHP/ogyvZxLbAnTKdklDlQOh4iyHQk4J07EMTyBDAHYxgBgbghc52d0w+UHEgY3gmROdSkYh+pATT5NoEJsCFXLwmZAIRYkHE0ZrTTUFabnKECoYiEIW9ho7vVGUgDigJSZBhjtgpmu0EYjwyVJAg3eiGM2KwTyoY750DCWgucEYFYGQgCA1kKQj50AmAfSgbU6MoVrNamhasj6MdoaQy6eWyaRHEEfWixD+eIc8h5EMgjP9gRxfV6MV/9LQjulACCzlliMDRFZ8C6cMYxhADHvBgDE1QZ0FCMAZfGI8KhkhBFgzAwKENJBZmbMVUB6KLymm1s0kBgFM82xEuZPQfLcgFJfZA2Y7oZyB1G8j9yjGCXLwRgcHIAxQK0gs6lGQBvbudBQvShz+Aoa0Cmcc8oMDbeAgkGQO5wigkAYx/MHUIwPjbav+BVu4YIhfAIIfk7iHa8ZI3KQ4SyAR4gUn6zSAXln3NGDYrTsFxFF3SMivb9lmQOZTkEf/AxTdiYKdc3POl/+zDKJyQ24Hk4R9X+McqPkIGcVRhCGSQRAoy+NTxdEIgQgsEdX4Rg1Q8Ik+hLS//ilPcogFol7IjaGB1cjpOSXxoBnWs1z/UMCd1yTYXTfgDOxa8EjsIQQm/cMcq3dGHbihWsCpZgPGMN4QMSzAQbwCSjIERjEAIbQRcPp4S7FAQaam4zCn2g4Pao8NJBRCLlvjHm/8xrlUOJBdtPtZK6QWEesUCBTFYgDvqihJWpIEV7+xGH9yxicHqYrMnccI/kOAOnobgH4wAHAO53AkqbHogQSDIAW8hYDOTukp7Yw4TCMKFIfDCEAbIBRU+DQwDiOMf4hgCMjoCMNtldiBAIGkPlPAPcPxjs8T+ByEzNOqORGMgPFjAYOEgZpI02K4RGIM7xrCAPzhBEoGbHQb///FpgshanJsVL+VqUep1v8cbDOLCaQtaNEukgBf1vvd0RRIEvhJmCuoCwusGQkhHr4bgHgQGX68YuAwIBKEzeMYudNEA8XZE3ey+eHSkMkPozKLhjHqNISwBjHEDriTptLWWGWW6KVTBnQIhNi4MXRpcCEQRF+brQAyQgRSIu5xR+AW2boQ5jBM9ogX4R8e5QIkfArETQRh5yXGOc4GoUhLq5GsVKjiE5hljaE+8BQuXXfB/2AC4JKfuPwxAz9k9wHpwsFzR4+7ZWXCBCz60wj/4YIkgqJ26BhgJPvlp9aI2gaYTrvUInkEOcPDA4MlRBOCe3pFvDy0Ku3h7tkg1dP+5cx6G7fOhGtprAMkbYNYiQexAOkgGJCe50gv4hRAe+guZJ6enhYA6zz0yO5qhIOid//0z6Z6ILgeD77PON9pLgnN38uDPm9hEBOyQiuyxgvbJmavpcx/Bku9+BChIA9w9EkLgkz9cF0AzL3JhBaENs/QG+Pt08/33kiDW0TQvNi7EbIf7K8cAQ8gAw4XE7qlAIPzC5Wxe+bHKtCXgR6jX+o1AEPDC+/0DL6SdSzRaQdAc/73EBrIEMKSA9p3dQFzX0KzQqIQfQdACA4KLIGQOmZHG0c0CL/DBEgiNJViC+9XarBVV8oGE5HVE471FB6bEuFHB6AkEyeUbGnQHEAX/QtBRDSKsoBTWRBEQRBG0RnLIYCwsQcFYggQe3/vNn/KVnIaIoA9yRxGNwBjAQT3AXbYQkvxMoRyyRBUehnLEYAdQShdKIBrwnfshX/h8WivUiwo8Q9Sg4EC8QPrMISOiRBHYIXPMQiLEghXMQCsclCEYzRfOXwV2hBmGSwMRTg+gwDdczgtFQSOmYkkMh3lwHCXoYSvwgiXczEFJ1lINxBd6xCf+SaxJ0NBMAQv03gEOxIJcFMYhoCr+iSTOABdeIh9gUQrMmgGkwN/B3wTuUtXEGqWoQQ4YQwQMo0AsSNxly4qUHzxUTA79QweUQDNaQsEEwb2JwzX2oBjuIhm+/4XjxYUl7B7NkAP4oWB9jCNBfEAytgon8MJQFAyl8AE8TqNDisR0fRpf5dt0xRkg1houceBAYENBfNrT0RNMLB3NqIAxGODlFCS7dcE/qGTFTAAbzGDBFFTe0ZtDUqMFfkRRTVet/UM4hEMVUIBAAOU/rMAWwMI/QJ5LLCBQrlH8ieAtisTUfUQw0IwajOITvhBBjBVKdhZLZs0LAIVCUooh2NsH1mRIzA0wiIM7CIEURADNvUNciIATdJsNiMOEHR4OpkScecSbjRzTjcAdfOMBQoIndMQI/NFWngT5NIS7ocQiJmZByCBHMeNC0iQ12uRIVIEQ4MI74MIpPEIzxP+FE6xAEtSAJtDDaf4DPdCDGTRPVJYEyYkgMMyi16nhEzZAKhTmP6QaIwnKHggEFmZOGkAmW3DBIcgbpQQDvYEgCE6jR8zf31HAJrwDdb5DaJYGPdQl1AEiSezlXhIEFUzl0JTkExLm0UmMC2hOYxInTBwdB8hgwXDhvDFnc94kQYihrW0BZ/5DBSRHdjaPR/YgbPpgEDBdLASCxFmOKnhCmw3EInYFMrLnqa0Eb8KFDJQa3cWCQs4nfT5kSIjDFryDP6hmcmAADsijQOAnTexe6ClB0C1oAVzAP8hoRyAie3ZEK86HNu2oitGdYCik4dAnc/6d9nWEOGDAKTSDHvz/w5KWxgrggOm5RRAEA/2oQSzogOXkZiVcwB7Q6I2yCo12KYq1ANJlAB8UTBnYWCeA4JRNWe4V6QjOVBM0Az0IhBmUxlwWAg9K6TaOQCy4aCrUwZZu6R60wpfahaEShDZtZSUwwCzsQy6EpSWyaQq4qfYR6T+gHqR90CaUximoBbGxnls0FpXSz4GiQxQQ6gVs6T9IwFWpRCkcqkg8ppcS5ywc5Jmm6aRWKq+iHgxVo6cJDRDNACHEQi7sgarmgqtqiay2Ra3a6q2q1wzoKpylwM5dq4oKBCGVz+hh0ggsQSxQQiKs6h506QWwwC7EQYQ2K0v85m+yZ91twyy8IrXS/9u1VmquhQt3ooRk/dAPdQIlUAKXXsAF9EDD5Ik4EgSLCQT4sKvDhsRvTgADbAMvzAATTKsl8sK1ZkAeZGRIrIrmNGWXFVTA7sETnOv3XU7CzsS7PmxialN7cEAGtMKZloCNWUIGDIE8rEI4iF1HrEg5zsgCvoQ8WkInjGwrtEAlxE/KWk4EyMEAlFYHtEAHeM1KBKTLquIS7AkXbAMl5OoMGKsXkYBAjJoUDETQzggP1IQYQmcQhIi/Jm2f/WMDQAIRZFTUCkTVEsQ1FIQGfAQDFIAxoAPwHUMRfEH5rcG2AEJJiAJNzMJLnmkrzAAftIK1Xto/OANI+Oyv/sNUcf+Z0LBALgQCOFjOCciBxGZUC0xABwxAHUSD5cQBHoAAAnjLPxzAAdyuQByAA/zDef5eFSYgHKzBcG7cW2jUrc6rJVJue2UA2f4D50aUTU7pyKqAGxjDGKCAH2gU97KuH7xu7OIB4oqCBoxDO7TDAfjAAWgA7/ou8BVB8DIgV5BEF8TqQIzDSnAI3SFdxU7umeZCCjCC8WhuZ/GcAfcrpQzNbJEWac3C6vrB92JeGuBBEXAB+bIv+6qvBrRD7/6DG/gCVmbteiTAOXblxFitQHDBj1YuZkWYthHE2f5DBDhD2sZF9JZhsxSUFSxBSvEBJfBCCwCxMK5BHNQCHiCAA4j/wjD4gPpqsAaYABcUwBNcwhOGRLNZzWKK8GpwATNYguRaYitkACjYAAF7xAxnrl2srYFoXwD+AwgGwewksNBMgQqMAB/0QCCgAArsAgioABfMQTzIwjDMgwaIgg/MwwG8QhQXAApYThue5ECUcdamiksEJ0skgOfIYCeAMc1aAj8wgqj+rCSvRfOV8gKo8YgVBOMdm0D05w3LRQC28UCkwN71jbB6Xb2UgyClIb4IBh/Y2SEELCVYgrh+wDMEgpH9AuY1wBrUg60RxCKwAYy0RDu4xwsKChugxDMOhAV4VDPRKI26qqpxgQP/aCu0wg+Dwj88VEFMCVyoMRuRwid8/4LHhgQYFARSygXq7fNAMBxiUSMcI89e1MsuV+kPzUAlFpSk2tg/bG3exUIVGMMz+MIv+IIccABaDIQpeATjdkQ6DgT7/kM1o+Sz/oMlU1SFqhrSXUDBTG4s8kODvTJckMJAkIIRDARS3nRH0DRpyLJHtLFPV+ANZlFMKjDNdNlCL7RAUArB/LKDaENGZzNIIK5IrC97LuoVnvQ3g0TdIV0LTG4wBEUuDAEJMMIoJAdPe4RNC8Qn/ANN6/Rq+HRB+GpHIlwQBCgO3rUh4E0wKGTNKiS1MnTBiC4vMAMzEATWksQS/61I/60o8AnFFME1J+BF3EXSGSdYYhYA0sGD+f+Wb8kFXAsEO3wCGIDBaLv1P5g2O/SCPNd0WrNDakdItgroLJeeOxbMmeK2xf6DMRZMLMQCOWsDEdQC43bFDRXEydJQ/L7H0f0ut1R2VMgFZAMxUFQuH2hsIVTbZ4eGHdjBPXzDN9iCQNx0N3yDeI0BcX2CEcC1ETjDiK7Dn8gyw+0DL6hXX+u2jeV33oVteyVCLoTMLrxBR1zobmoTY4fPcrsHwVLMicyFsSaCL88Azm4DMjgXEpAGR/7DNziDDdzzUf7XO/jXI/jDAoi3E3TDf/2Df81I2woEGxfEPvyDPDQcFcyAMTAvQy/1hlLu1+7FDuyACshALlxAjO4BJcz/wTAcuBazBRFMzAsEM+VKVWGL8T8AVWk8AnijOFL+QYZnuHLIQxaARhbM+D/ItyVwR187yzYzL0GgMyX8dglcQCsQbCUkQkf4gJIv+UvY+cRYAC98beVSwj5kQHajMWnA5SNggw3ctC2AQXk780CsOEFI+luEeZgnRyzLeNplIuUSzFKfqTQNRCtUwg0qLZnSwSskQxeIwjz8Q57rOVYBwAhQQqRilrVmQSE410DEcEjQ8CivBFwKxP2FgxnYQAhgA6X/w4hmzqV3RAbMuDxQYyfIGH4bpuF44f+tQh7g7z/EqgeM1xIJCmJyC0PEAoQLhsZmAVlXm8CNxiOIVz34/1ewa84ajUQAZsGzA6C93SA97d0NgmDO5uwqgIIsuPqrU1RGPESDy2rw7MAhuFcsTBC+F8LzXvhAyHRB4nuZ4zvHZ0DHc/z/efwqxANzCcTf2i9JRDMnpGf4TGiKecEyTBRo7IIAqEDAbgcvgHkWZAG7D8R2b2WzD4TG/8POF73HD4G6AyA/aEMGQMMwlIIGRP04FHIHw5CaiYTLO6vEGBNp7AJDqIB/K6fHHwGu9Txz3B9cevlbkDmZ00Tbt8URaPo/dBCZF/02ZMA28MMqDAElPEElOP0FR30h/8MhiARk/wMlh49myDxbaFNJa86FtAUe6FAuSBUAFj0yYC6zC/9E3Gt60LdEG8AEP4gBPxCEpXd+Qdz9jPND3qdfLDxBAeTCE3QAkkN91EN9KZh9VmX9xUV+WwAAzffA16KBtYJ5IWT3g4nP24vBauQaP+i93kPAKki/9Ov9Klz/HFy/NlBsRFvZG7yBCpSA7A95B6zCMAT+P3B7Z2Wxy06+ADAEC3xtMBR/FmwDrucBpGkO6g8E8wPEP4EDCf5DVhBhG4QLFx75JwYCCQjbgj0LdDFQLC7bOG1E0BGHsR1vRpZ8Y6HEhSeVLrSYI6qLQFEy/41geBNnTp07efb0+RPowidBiRY16tPc0YUMBCYSiCeAgH9uEvHplCFLVnnyChXK82//jFKxY8niPCjwrNgsaB3yQ7YKVIpgO1TA4MJlEQNODPgycGPhyxtMb0ieLJHrSYELXEz8K3XzzT8AZSlXtjwWBpOhlzl37ozn3643I3gZM8RLHtYs8rIcWesZduyCEAgeTDtWzD/atPn9W7Vqm7Zt27gwQMDgrhsQg0kG/mKBhcoCAhsXdCBwx8DJsrl3F2vhXyzv44Gi+udCKYJ/TAW+EBDImJ9cfAxlyMB6W5ZCrf+9Jv//J4XMqgyZ3JBBppAhUiiEn1X+mQMuB7dBjguRmCPsjcmia+WJC2ZJJ56YZvrnlQT+iUygXSQDkEWl0mgRxhhvmoCLf7gY4jhmNuKC/xdDgrFkn/uyykIMfvjhT6CvZISxjdwEaoM22Rwy6Ml/2jgiA154sUTLfeRpkI7feMEuMpJ2COSfXHJJhBdtftuGGV7E2eaVV5a8E8889dxJrzmg4WSIf4bgIgX78stKDIjEyGCIrLb5p5CFFthTttwEJG9KhdpQyMghDKDCklwoySVULbVsgRdUTaWEF0pcpaSV+QzJRRs7Kb0V11xh3GaOOcL8bRUIIHhrmyFGNSSFf1jT9b9LWUQmStv+4acNfuTZshNKsnU1224p2QPWXFqBtZNxWxFnlXiYXZfddjkbQJxn3lCBFy5aubcVPlqxhDXW9ptyoCbcJS/KzpwteP8gCICTJwUDROVWW1glbqXccLlQcjzQBt6YY+5qjIWQfSgxhA80+LBKtdZUcw3gjjlDhoSYddttPIQF2g0CI7fK4J8UUtBS22wp5sVBhJ6JbZcvdpFqJxRcfppjC3JQ4Z8eFvKDC3EQYGYbIkQt1xBKgsxqv36RLEgIo2yAuqCYQSFBN4liLPiKmaE9UIxtLOnEkCp8myOPBLow0TsVe1IBBKfZdldxXRt5SoXIR5Cgpn+q+afeIYbTZpZWWw0aNXlcy0JI/yJdKCxmpRAIicuiJAEUOkCJm+badUu4M4SdxXxvVtngYoABgB9AV8MNXxz5PFVA1Q9eZrmLl324yHL/CC25tCTUQvlJ9IgjRM8iP4H8e7r11juD+x8SZH87ZvQJTv/maflJYW9LMhC5AE5emSMBwZlFMXkBVAoLlAKIfwgAANUgjZrqZb0tjalL+zBSzqqFjCOIoXui689rTicQebAoAgOZ1KR4Uj6g9IYgu8tJ7GTXvhatAhn8qF4u7pKLEdwhFh9AQP8KIgKBgECAQRTiP+4QFAP+44gAAMAbPsAjrglLIsGSorCoOKwmnWVKkdKiQI6AIGV1MCfOGAgFBoZCKgGFNiyUHSNkxoiy1I0gRYvfETQ3BHEY4w0CeEMUYnGHXHBiIIQriFQIOURDcoyAZEngP6JwiFD85gpQ/7yCREgQySraRiFnORtEhtUVgYAxgKCU1m2AAjs60OEfoMgDKGa3EJvxBI4DeVOx/PCBQOABDwLAZWTuUESdCMAXUgnAIYnZLl+SpRqYyM4/UIADuFzhN5SMCLSEdZaDoHAbyIDmNpyAAyeQoSuF2MYRuqKkTUDtBv/w4RVIScqfzK6VAmFhPv4xD59kkiAQqJuD4KLKKxRLHFEQQAB2EQBfGPQfIHjBHaz2ywMajmnFjJEAjkeQhvaECIdgVxSQ9gyt9YoOvlpFAiAZrEoC6x/boIYrNlEBKUihGas7RwU0IYxMuIMCN3AjCS1TA8q07B+xZCVwgOWW+PlEjj6J3f8/8nHKU7JSlRECBbBIECEHhWIbCBAHEQggBwIQIBAH/YdBh/nDn1zCF6GR6JLQOhA0HeWYueJo1S5TVgIURBxfxUIVCEEIT5wBBYF4wRmUQAEMIKEZ51iIYl3q0nA4gTyw0Ek/GNK9MwrEUnS4QhV2UYVtMOIK7JxZUNynk1aSIA+oFUixqmCRN+wCBBSNikGj8NWvEuEfd6UACIIp1gBcYq0CfIFAqAaUD7TrDP8obnItU4cPfOCu/ziuQICr1n9UVyCGFUIzxPiPZjTjH+dIrB5WAItByEiyRWknKK6wC/fughBXeBu0oJlPnJTWJ3BjZfug+k9xVCEKIAhAACL/EYAzPPcffhNIFarAW+BG1Lr/EEdwO4bdnxCCIGRs11u5M92FXAIFX3BaHSigicT+o7vh/Qc9anBenJgPKD5diE9lLJAaM8QVQYVUQ6SVz4OAQhy+cO9BySGOK8xhqpU0LU9Y+Q8lwZN9EYlIJLfpChREQiBn0LDfjvsBBRckrT6xMIXZVQsyH+VxRinsCn7wXe+C9xz0WMF5XVyZ9P4DFjWoAT3ooQc9hFcPNUhCTlzhimcM4Qr8ACMWB7LeVVTBoBSVdCA8uo3fQPUf61tFHp7aZPjlYQ6pLMjsUAu39sUsD3BBxhA8obE0l7UgHkaIxnoy5jPfeoiNAMQRgaKE/38owRMrrgB3B0IP89b5HzkeS573rIdzKBYhzfiBd9fx5xqsAM8DGcRKmbmLCdMmLaSM0qVg9mhf+AKtAaDBP5gLxEAANhC7IEcVbiAOMogDB/gmAAWewWACzAmOp4zHK+JxShGIwI7PCPAbqkvggWD5HxhGCBbGAut/hBnXGWcIrxFi5iWlWSloctoNVjBsxTajAnrGc3kHsQJq/IMa3AYKLJJAjwpA27v/mHZO2twMPdBDINh2BTU0LBCPPmhYtXEnWgRCgjkMYWm+oIHizoCmFygBuMOk+D8wIN2IH62saYWvQHAwEPXgBNZphjgWtv6Ptg/E1kXxuMbpThCOF//kcdkIIgoosAI9VGDYAlndQCqwghxnws88wbZAhCGQ74J3IG4uCHghP23w7twZcfZpPyigg4GEQSAYIIAHCnKbgxzsLex9Bgp0MAbWs/sfw73uP0AP+oFQ3Glx5wkKKnqTtwvEzMDVfd3J8qIXDXHugIgDICCOEAPeHXlkFAbgiT0QPYRjBUnAuUC2X5A7o5ggkAdKd3cuEGc0w/BF/0cd/nG0gdwAByIQJEPgOCyFoVIchEWB7P8xd9rffv0aZyGUTSDSiQB8rSD8j/gWECfCQBD+4QHFohhADokWQgGDCANcoQYA7+SaQRhcwe/MjycqIDbOQYwqoOV+bd0Ggv3/6qDt0ukfyMAJPEABVkEEVgG03CaV4EY4hgAHLGL/UAAFLuESysr2BIL9mIsgMG4A1Y8BnxAoIhAKc6IYLvAftqDQqK8CsDAJxC+MZKO7IK8C1mEFMoECtsAoiuEfimHAAoAN2RCtnMbzEILDIJAoYHAFpxAhIIEsBAEBBcjXBFAPCwIRasEKBcIMMCATXC4TSBD8HC8num8gGEsstm+mMmEQyHDxaEAJpJAgCBAnakENL64KBYIG5hBt9IQWgmgVKQPG/iEPkUcI/lApKPDW0PAfzKAfGpEEvfALxSLFJJEgerHwVuAcBm0g0gYhFg8ofgEWn5EGYhEVYwQB9U6A/9BBFZIHDtoFHQoC+pTCF05A6mIRNjxvGgeiFhBhDjnRFZxgBRpPT7qPsYRhBbBtHW5CEzwRV04gRlqRIEZxEIliDQRiIHMlG61xILqRLMzsF1aQHGEDEf7hGm4iIrfADDKBz9qlGZJgEJJAChzxH/gxIHmiGPwRIcUCELLhcaxhJHNiIrkjG1LyiFiyMpyRIGyyM6whIkPyJlQhAkbBDP4hCQbtnNqlHgdCGAZBCHZSB14xE3CRINwBIbLxH/TuG8kD+nByIXZNKVRB71jyEH8iLIWoAQTSJ1IBQBTyadCyJ2kgHMIhEwYN6AZGGO5RINahxARCGRFCH3tyIbSyO//iIA7+YTB3ohGsARBe8ipzwhqyIRuo0jLQ4RqsUS1xgiYJ05DWYBv/4fgGgi0hky1bkihGAQfCIQlu7GlIEAMQ4QR4qiD6Mldo4SUxkye4QSAg8ye60RpUISUj8x8UcjZzAjd1pSyJYjM5kyDQUhWosjO9ozCRs2OacyA6E7KwbdAyQVfsEiEc8R6xcy8HYvA6pjJ3wjZtkzZzMxsUEhst4yUlUyeocjCf8yb8MXnkUyBwQTRvIhqm8x+k4R/s4B/YQSAU4R+wkyf0AB5xZdBWgA//QQdE8mnA4T8WkyESdCfU8iSPIoQEokHz8yY6VIimAQ72kyDFiEAHwgyQEWr//qzxaqAfVmoLwtNDjQLGXvEmFLMsOjQVKDTjTmEnTmHaQFSApmEg1qABHusPBOIP1qZAjUI7uQMkGWIdukERkkEE+mEFzMAVmiEVXPMfvBRX7JNSXMonuvEaglMp+JAH/iEVxBQo/EEggPQffJRj/PMf8JMnfHRNM1MgeEARwEBJUZQnkmAdCrWlCO8eLVQoL+NJC2IdBi0c2CEfSIEReoERzKAGMsEMSu4RUywgdWEgWMEyRBUtQxMn0BJUlWIBpABMb8JH6bRj/FMaWIFEF7AB1sEJkvQfdFUguqFJF8JX/2EFGIFYPwEMwiEEhrJQEbQC6pLxyoIesY0eCHUuj+HRV20gGSZVIHohGdjhRYdSU1cACSLAFwcxVTlDVDkzXcdjQ3UCP9+BSDkGP+2gVm21GwA1BApiU3PCV5OgSknhH0gBYP8hGRgBDMzAFlagG7pBRW9CUXeCI4dOKBvvHu0yKAlWIKCgF9jBDF7uRQVtEakhE6SNTfVEOgGEFeTzXCkjDlL1ZBfiZY3CHwICACH5BAUKAP8ALAAAAADoARkBQAj/AP8JHEiwoMGDCBMmFCBAYcE1A6dJ0+GwosWLGDNq3Mixo8ePIEMSxPOPpEE5AjuIXMmypcuXMGPKnEmz5sxiNjc2yMmzp8+Kpv6x+Um0qNGYDQdaYYkC3a8FNMacMdZjxBQVO3ZUe7P1XzUAmDC92WEBRKBAzz5w4RJKQZ6jcD0yiFvzF0EmdP+lycu370A3Au1xVCdwgMhJK5UZVCxQgl+QDh5LfpxqIMSK14zuFAhoMsbNChNldPwvFBs3Fv6V86JxUjXEAf55YVwQU7WBrBOWQ3hM4G7fBJcJBDAlV2mBnDy75PCPw1zl0Duiu9zyHs9aAztHD4nO4JMRHKeU/yvXW6BwhADSLz6fkH1w37n/HfstMP72+/jz61duvaOqAG/0EMsOqv3zQEXgoWFMIAUqc+BLyygTYYH/LPObhbMVRJtXBTUUSSQCEcLJIjUxt9+JKFoUm0MfxBTHZqA9Zl1/HKHwTw8aTQGeGqptiJGPu9GHkI8CTfGPkRw9CMA/b3xwQwQxJoTXdhwwF1SKWNJEY5Ys1fPPNBmhVJAKG+VQ5I++jaCCMuXcJhAat1BhyAjj/abYFA8ypmMsVPxjiSGBlDMCeA8gSdCDFFKICQDPoEAdQfY8KgOXHSWgAaWYZtrlP14OhCNBfvwTKkE2FsnjFFPw6BCRBwUzxD/igP8n3giG/FMFGgL1SQUwkvxzCwbGGLnbA+AZwscIAAQSTK1UoCHJq7dIAkyz/6AxRCH/DBFMRQd6EUhTcIQb7hprfFOupuime180+VUi0CwtUALePzzOW+QIx9Kr70bGDBTCP3300YSv/1BBxRCS9DrQGAtgw8MC/RZURbXPDnHLLf/8C3AfY0RrAMIDNSHtQH0CYxVB5RgZSye1DmTMLd0N9Ii6ND+Gi6YNwAEIiHlFaRAXAk3wDy8zqPpPK7UGEwwOBC1I6z9BXJRPR6zogosdVT9sEMYDjYPQFQRhIxAFQwzxhyIGUNFJMKj+A14QlFQLXix0/2NMFOSM4Y4/j+b/ZyJLB9Qs+OAYcTFLLiMspUYwQRgQBDCW/AMMMAg1oQhBfUpORTCDukywX6zw4I4TIw/0uAEZGGAAMBlksI07umzmJY324ET47bjnbtEslMwAXicpqP5PCh9dccQ/TcQQw8PL68LDP+CAY7VfGQBjgDwpABM1yYMaM8Ya9cD4z07kq1LzHv+gj77u7NO0Ylyx8PHEP4nwcmwrlqTAi+oGZDv8R5SriB0EwoqQFDAkmTNIEOQUCBXwIQxraEADrEM+gkBCIdlonwZ/wocyTGqDHuHDPyixDz7MoBMDGUEw8vcx4v2PeC7cYLMGxQcs2EGCEgRhTgKXEMHo8IcrkUEu/3hBtBLMwIgl+EcuUjAEJmYrhhZZnTiAYQNxUAADNcgiPQQiDJv0z3GmC+NGghCEQakhFs8ABw5z+A8fVoYgPCLTP7TTlw0IhWk044Y3BjclILbjIiiYFB9IyAcjtmIGAslfBlKQgYG86lUGcaE4JCEIXLyjGefY4k80KZAamEEcwlsJMNAwKBW4gRw3jCAb/3HAgVxgfhd5DhBdcgkqcWR9s9wIDJbwDybEy5AzECHwMjCE1mFJeTHpXxlHoAY+ECIVE8ThPXRxhgK4SyDXzKU2t0mUKPyjDP8oQSsS0YIZlMGcM1jWPjKQBWOC5Hk0U+acfHcIcsBhgnE4wxMqUf8JSuzhmrt4IzclUwTB/U2bJXCDH4h2yEMCr53yyMLxWuKPgYiNS48c3uaOyIcWJIIS/QxpLN4ATQkuQA4HHUgYBto+TgzFIbDEJkvgARI5QqcSMR0IFziwjxm0gg9ARV0h2JmFK+QhHAsQSAUE4gyDNPUfMYiAR2IA1YNoTCALGMNTx+CQq9IEksPbRwqCEIxWrJCIuTBELtZSJTbMggOzmIUflKDKOATAAlwYRjw0oAEojOMAf/XBK/xwCEoQwhe/eMovpKcLONzwpAYZyg0+4gOavQBFb0gXexDTCJmshXc/bUUrGFmILJT2HxDIiy3+8Acw/OMTArFFDJzhjHX/2OK1rhUIKf6wAhuYIS9ZaOfwUgeMTqAhnb4LxKBGkM4RoKETluDF8MCahX8MtZ3byIA8MiBWA7CMD9tqxT9MSF5DiKMKVTCGMVTAIIKI8B/QYKlI7PiPRbxUvjnhAjN4kQvwooGd25CoPP5RXUbUBBs3cwg2nGEGMIDhD+t4xDv+UdF/THhmApkw+7B1vOCW1sPBzUJE20li17luG/zgxz5ykYsCcCEdB9BAOyorEFFYJChBcYFPQJAaoiAGJgX4h7uCrKnMHmQZ5fkILLN5kBe8QAUsGOIM0GCJdZb2tARxB343IgZkDEQM/wCzRtpAgm1U4Sw7CIRW0ryDWAyA/xMMGBEnOADnQ1jAAll5A553oIInXKDFIIWGLMYhCg2IYhwOsLFFSGRfj4BgIAS6SHuNwrPtlIJw772AkAUiGoEgwJFDs18uSJiBD0vUulsuyhHaAAFQgGIedADFP7bBC2BELBb/eM42cs0GZohjiLyYBS/2wQtKtCIXouWDaEXbiVYAYxXziIwHBGJkNxmERLpb0n4UXTMYFCQWXNAGL8Qx7H0wQx6rSPE2jmDaf3TY3VkI8ECqKxAtOzXVM0ntP1YBAQi0gd8QQMYqWI0MCHSZH21AOD+QcQR+HOEIYtgGJeTEhTnMowulSHRk/hFpfHs8JAT4RzEakcHOgOUfKv/oAQv8XL99cGEf0SWiJaLLjC4LPMUPbze26E2QiQpEYfhBgkxIIJB+p1bfeUE6aonOb36Ig+a8eIIbJjCHLiSgC0QBgZFRJI1/6OLjHmHaB2KjnWxEogriEMcQ1o0MfgAcAiSI+ypIAPe6I70N/2iDmAfSb3f7vBBe3g8SkqoQrrYEFPmgQ6x7EfeBGFggRIe8ReiuEVDEehueAMEudoEHzu/i0QNJDthjYpKCfOoMeKBBzZ7Rgx684AwiwQMA3tCQXdxgGx6YQx7mkA7dh+IK4rhBel+wC0Ks4go3qMA5nHEOgjTDGRVIQiZWEA4nbOMKXejHQIR+lBUMZBAYQQb/CeigABGALRR5CDhq+T4TWQskHvFIgAi2QYAzeEIFUXgBCBgSgABEov8BIADk8A9EUBAFSBC+IBBJIRMUwCUh9w+E0BFpAAjvoyIKAXrYcRAPSAgPOHoJKBC1RANKIAg2gAEVcILM9w8V0FR6QBCuMBDa9w8i4DX/8IIbUQOdJBDroAfN0AwE8QP/0Ax6QA9ZVBDeBwv/cAPksHlVcAWrsAr/EHh7t34CgXd5IA67EAC7AIL/kIAoQAFk4IR5YHkkkAckwAhzR3RlSAKgoIb/AApjaIZxCIdwWIZ1aIb/wIZwtwp0sAoecF6B4AuVdhBKIAAfOHoeESl70R10pBDW/1BpKKAE/yCJBEEDiKAQK7VSlPgRnTUQ6NCIFTg4FOAKmXCC/7AOAiEFwuB93aAHS3UOLaiCBJEENbACKzAISDgQFdAMS1UQ0HcQT1UQy3cQUvAPONiAqlcQYYAFBIEDN+CMOHB91wc2q2CGaDiGr4ADZxCJ/3AGl0UQkhgGGDAQGMCMDsE06IhHdfAPlwV7/9B/AzGIFYETtoOIBQEHGLEXeSEIIhEzcfAP/9iIOUF4MlFLBnEDTuAKXWQQzecZ4Dc2/3CJ/8CPGUELCpGMA4GRGLkRDXgQG7mRP2GR2FGPkiGR/2B4A5GBFiEE/zB4MeEzaxAuXzc4GSQQiCBVAv+BkyChj/8wQBehC2mgC3GADitADTiYBBvRRV20Cb24EqhYEU95ETpAkBuhChlUkyGhCibpEsWYih7nD0CYS2EpE9egCtzwD2VJFw0QA05wOTAoEN1gEHGpHwsZlziYDDZYEE2JKc9zCjoJE5kxOBg2EN+AInAwM9/ALtzUAJvgBLc1EGYQDjiIgxWxAuxQEMnwD4xACp9ACppJCr+1kCxRi9TwDysgDEg5EMLgSZgJBcngBLaYBK5ADadZA9JXlCugB6dgEfrok+1zljmhmAnRdf9QmAPBk+rSN9/4D0Bgj87ZEkLznNLpnAvYEiHnMx4hnAhRnfiVUog4F7KUjxj/wZ3TyRdPwAdrMhDlMAmrsRK3sRvxcRU3UgJLYC+PEZ3lmUvGWZz52RGhoA0CkWQXwRoEKhu4YW0HYR8G0Z4BqhDVYCSdhiVY158+YT4C0TcG8QXk2RObsQYCaZD4gZ0HEaEIYZAjUAJP0JwgUQ3HgAn/4KKrgaAD4SZeIKMogxDnISQI8WNvkAvJoWO4450U6hAWeiIgYg0CIY/QsSUakUEkkVk4oqMJYSjg8RtBEhIWop5e0CZf8Q+z56UCsSKHWHsDsQtJ0RACEIBR8Gljo50vwQETIKRDKjgrsp8GgQelZ49w8B+xUKUXkTI3aqUDcSDuARJXyhFSWg4uOhAC/0AIXEAAqYChc5oiCaBNIioZJ7CcCDEq/6AKEbMR4KEMzWkoGlENtpEy8YM4GTEegWAMbCMQtMEqA0EbB7IkFkAIJ0AzVzKpRwERdjpLXtIpDQCS/3AIxhGBFWE0CaEYhYIoCIFrhyIQc8IghoAGE1MFCZNe9HEggsIHxjAeAvGpaEAF5zUDhjAnO2AM+WMReCIQ3zKTBbETYDIzScSr9ppLSZQI+aICJ2MQPFIvpAoStxAwt8A2KiQQE2MrHyMQpMMxz0AggvImfcIsBWMAijAwGdMHCVMtwJACvXJbVWA0UxALM4AkjDEeg9ImXjFp0HOv0DGhKzGYLrsRifAElP9ACWZSEFrGIMy1EWBTEFCQEJIwBs9jB7jwDQtACFXALP2jCH+AsQPhBGBwBa4lCYoABo8nEL2APDEgMv/QPylQrWqgrP/AOVRgHBODAVQ1s2xLEzsxgWGqluPjEGvBCypkCblgrpGTSAeRsHsrJ/ZJELfgC3rDMBpxM1YTA6MwCt2wAGuLNQKRYBURDv8QDpuwCQvwMDagPWuzA1OwLRWbAQuUK7YCDOJADrEzt/vBHHLatq6bEUAjL75jCJYgPAGUEUZgEL3yKqYbDGj0D+SwWH3hBMETNVSAOgWzPZxjDELQAOEjEBVUQcz5utSrLrEgA1NCCS3AAjMwA7UbPFD/BBId2UqR6xKS6xGFQAXs1j8KZCvKFQvkgEOFCRGXKhBG0wj4WL36eyJR4AeJ0L3RZQDghUIfE0q51Cxj+0CqRCP1u78usQwFtR19hIgtQDTdm0QlAB68EDxNRBBgBVYFcbsGwb4Dcbs+BxM/yxJUsFxVQAMRdA+rNBAC5cA03Bd/ZBEoAAPi1ALlRF6I5CdM5EQgfBDEszoEgAT+IGEUdg47KBCxaIQiAQYL2YJbRISfRMIgETVzogYjgEaxs0aqu5s1bBBIqh8mInou621KtA+tQLKtUAIipEjFVEwX0T/iEAJIQA9ESA+p+RMvOAhkAHQegcWSwzmDgkZ2oEoN/xBB/3C+Y7wS7OGmdNEKuGSP9BlOlGA/wbTJaMALrfPJKGIHPpiTMPEqKzwoufAMN4RD1FQAIPXI+KYSstoSTFYTN3wR4CRCxWZE52RWqNM6WTDELCE2MosiBhA8luA7+EIAYxAHSmCz/HQB/DRSJVURivlGn3YpsDwTu2oROBJktSw4CtoSsXAInMALbpxOubBO7QR4G+EMa9sRVPWX+pECm6NC6/xyiZALKPAiMCwEA8AAAv1WEzABfnAGdbUiwyAK7dAOBxA4N+wA+AkHfSOvazCWuRoSN3zLFNrNCAEe4VwQLGsRr2ACJvAPNEVTCsGpAtFjH7Qfc7FreXtIVP/WOgF2BIWQB04gEChZE7BFEJyZuwjhmcrRSCnQbCrUCs12LMqcA8z01FfBxcxlBTPAAtA6EIiEa1ctQuIlQoaUCOamDfdVEKA3EHGzzW0bV0AjbMFUBoaQAqUVYFjWExVmEAkWDrn1D7JFEBP2DY9gB3WdFwOGLTs3EMQkEJC0sB6MEBIVXAQWXKUG2ddlYsQkVvpjADO3K5YAOSnASGuXAavwCtoMEvE1nUSGLtXAEAQxzitxTROca//ABQwwAftwCPFDBXAtD0cgD9iCahchVfEsE4FNEI4MHXgHZifsEfwgENvQdk8ICk/Ih3MA3emwCttgCWc2AllBFn32T9L/XABsIAuXMtr30WM5saEzqwD/oN4swQFA4wa8wGzALGKnJhBgYwM1zHPb4M5tV3AkkG4ZIA7BkAvGUAVcwAnbMGcKzgC5QBZ5pnV6Ztb7MAvERgl8YCyc8AqiMAfQ8WhlXRPoHR2X9g8bVzNPsE9xdQi8oOBCQeF4e66GwE4RxW7BdTy9bRBUWcM+R3AqljoGcLO5QAVAbgmdcLNGvgeUUOR70GzIhmzGYgmCJgsCIQtgtYXbFIpti8aN8CEIMSk5FdvMIG7FltnSpduNDWKEPWAWkeOPweYroW9IF3kGoXQigXcDIeeRZ3T9NnD+5m9tgAwJx3BDQAlrpQ0K8Aoa/94FotAF8bDeRdFx22EH+YucF2ESVl4QgDFQjdAINEABVYAvQMUHuVDkmZzJwDAEXIBidLfq/cZqbYB3dv5u7kYQ1aXmWLIJCMGS9cYRiCdrcSfnfrEKxPSob6BnPQADbvAEDLAKoTBtBqGpaD1QgJAUxrANJHAFfQ53kfd4UIgQyFBwoBB4s3YE6/ZwA5HcAsF9XDKXGuGGCeF+7icQ+ZAHb2EQ9V50BgGF/z2G1u0B24AAA4ADcnADciAHBEAOnXcQ3hTtCc+OCz8QI62BWPIpLgGACEEByLgLWIAD0e2EV2ADwrCC5/B8uigQ55AEuZgQ6m4RDwkSLU8Q3R6FYf+G7lHoZbt3BVhw6eJgVE/YdwQB7Hn4hgextfduEFsrEK8wEH2IALkQBSCAAmn6f/9HEBGYsP/QIttZEGLyEZN1gOOYJR35D7quEZReEbVw9iRpE3iEEPX4iScikBzpCkggmusAC64wCHif90XpCitAD97nEA+JhIOAg0/8Az0YhBrRVOeAmn8/EAmIAYRAAYSAARRQCNWodPy2dEq/DeTgC5tHA76gBEpwBixbKmcg+WHfgGGgerGRgQ04bTu909OGADeAAZ5ADgwSCB/+D3uU9rBMI/DaEQSpehapEOvIEiQJCHDfEj3tEAsACP9IE8lYBzfgCnxcATXgCq7QlA3/+Q/dL4sWEYwKwXzQl4IDMcq+SBCZ4PgqtY4rdfH/gAEZnRBj3/yHaBDkkIwZqJICARA3/rn6V9BgQRQoDDY6COjgw4O+/kmkBdHiRYwZNW7k2NHjR5AhRY4UGcdgGpIHf6VkufGXEFeukmRK8k9YS5bnQHazeVAHDYNClAjJtNGaRqArcS5lurFYU6gFwT0EWhARSGcVInRsoHGNx2lMt0ZNmcqg2YJKC55a+rUjKzgF/7BTpMhMjX81eJLle/FmwZtbCi74p+OgEIOaLKqyOPXfL8Yhs/2LvPRaX8yZU7I6xaqgP819eegqiMuO59AjUac+uGaTkz+2bBXsF27v/8ZuK7rx3PSvd82HvT0C3yjsZpK//2oSTxKOkcFeUJyYMbMiyQpX4Sr8kwKS9EWzPAxCYl2+PDfz6Q0K4Oj2YDT18eXPp78UQMHvB/38m1Df/38AoSoiQAILNDCqHAz6QiNC/mnwQAgjlHBCCiu08EIMM9Rww3sM6rAlTJgiQocGulrjw39GkGCEgnbYZZd/LPhnBxBeLEYXOOD4igARIErAwQ3V4wKBIIuMyj0jM0Mxo0MMqgezAmIZIZBqqgHgPou8yLIgTLT8x4tJqvkHkylGgIEXLrb5J4AkNeOizY9k8C+SkI6C886RgHhoEi81EpOpcsr8p4SCWIywPzwTpf9wSUVxQnKjrv5ZbaM5FAhFnH+UMWgSj/rciNOCOAUVonIymkRTgw5p0kgTGnVVyX8efZXAOf7R5oMdvCgVpDD/A4KPfxI5yIVZi7XQoYJktegy+pTFU9iCVu1oFiICmWTXkDg95sov/9GW1FBbKhXbg8QEQIU3/+HEWIg4YLfASEHqMA6GCmKTtafofBejHJ5g0dOUdj2mmmNQ/QdbcjVK+CCEMfoTgFwY2LfARRb5h9iJ/4mXI5PsfciezPLNuCD2CuJDjSkyzfQBjFguaIYRPGXZ5UkwuZJbLkfq8xiDGj54mX8KPvggLP8ZYN2DnrwTAYv/SXdkqFvS9x86p5b/kFGSxBxhYYtKTbkgY0p9oByAl/JCmbF5/qeaMG/+B+eH7i0IEHQMMimNOMgh8h8Covb7zvz+xkmVAECIJRCOUNXzIJaXKQfogiCHqmyNXO75IIP/AWGApgX3HKJQ/iv5IlU8+bylyWIZaQbEGbb8cote7yhzg2j3aBnaVfDjBvJeRfp0j35UAPhkJVSaIywMIkf1kEaYoSXJy1GBBUM1yjzQEcL+OqUe+t74TlOITxTr0Jyl73iDJMgs0BxU8Ijrt2Hc4flgDOEDcU0Xt2iKcgINBo0gPK8gtstIOSyHCWPQwHwbCp/42vSoF3wOfR45wUb0BxFNPWAKssOgCoCg/ydNpSwYhhoBsFqBhmAAAxjB+MfXygEEDf5Dddj63z/QQAUqGOMfwWjFCDQ4g2Ck7IK1M4jLAkGDb2jMIk/ChQOd+ETNPOlJJfqIEnT4DzVgsYWzK2DXpmAMNBiChQdBgwqrcItg9K8gGmSRIQIhAADswBAGqQIahjAESeAQDSkKQkGo4JFJBGIXcGjAPUpUSCVCUZGLjIoUE/mQfTitBbPgBS9UFQspHQRlWeSI5Th4xX80IYiBmkEnDEKFG1ZhCE24RR9ugcY1lqkV/6jCCEpokBum4AoFucIVJFGQKkhiCKGURC7WeJDtDa0cgRjBDnYQiDeA4A3/CEQwlJBElP8wUpt3qoyECkBJYLnPChgpwQw4acGu/UOA/+iDK6tQTUNU4R+oHOZB+jCGGOjAGFMo0xxxico/rtIgQwADGAqBRyqs8pUWiQUvZvA1l/UPk7aEiFr+gYdtZlSjTJkAF7iQCxZo8SC5wEEVtjcF92HkCRCZoyL+8I8QhOAWNyyIQNn5j1t0YxTg0IUdeKCEYBjjjzbE4R0lcYuDhKCdY+BBDG4xzCYYpA+0/OU/+siLIKZsCo4o1BQMQQV5GmQMG3VVF54YlwxJzKO8sKUanEeJHv7DBv/gwfKmoIYZUAFYGpEnFSSRjI+E4B92KM03FrAFChCiCYtFKkYYQQKMzOb/IAYoRApwGMRztoIKweCDJaiQAmCMQUffI2tpK1QiOADCGwAiLUQ8arIRqCEWlDDECILRCQP8UU3/IEcT5BmMP+IwRRYJRhUw8AcwkOCgIWGFLlgxFXcc5DYicYdMW0kGYPwxGDvg5z/8mQIbznKMVQjGLaowhjW01rTrLVC9LsQAXkjJeYbghUHk8REqdMISwXhed/+hglhUQSIQSeI/mkjYizRXF86VFGmaaGBJHSQcEjYIYXlwYZ8uwAZ5tGH1/mGADOQ2u2AdgjiEkN5/JDEs5GNvizV6gX8woAW2ZNEMLAGMeV4Exzo+SD1XGIwsqqG8Uw2QeK6ARz/OMwX3/83AMIPxDNHaowGOLEhY/lELF2fZtLw42QxszAsDGOAfOyZJE8Yw1qhW9xaLFQcFmvALOyD4PwYIQhCWTOcg5JYKtjTGGA5ZkHgprZuzkpOWMyY3+tzBIK2oBBf4ADP6GkAc4B0zS6C8iQUXRDwQLk2BspAFMZ+yj24cQSyEMGUqLsYiqGIIyAwNJ/W+OiOVaAEl5puCMIea0mTZNC42TVf/VNUiODZEmdxADlTHetUHYbGsnT2rFjh0BPTFNQrFHOZh7lpwqHTrE8iRXip2RdkFGeKzzT0rTD6hAH7gQyxmuV/bmjLMwg0zeLU9ss26lQ/PAHdXQLaxVJju3AOPWv8LWjCDcj6vBLb9B67vfbrajoAFVfjFNwo5ZYJn/G8ykEEuKolwhBuqE7wYQgrAW0+RCPsf4hgmDh7i8rlGBRn/UPlB+rgRHOd8zHuOLSE8oYtDusfVD1lphDZwsQa6Shoax9ALZFCCC0R7Bo9eOKFGXvKHW8TevzRACigQAiRspRnNKIge/kEPsiSDHQOxgQ3MQAYckAG7dF5KAGM7gg+c+JBUdDVaDEKohyzQPBs4uimepig7Md1CMPhHK6T+aKr/wxIpyEAKUL4RAwBDHFI4xTv88Q496AHtmkH76A9SAzOIg+4FsQRJWr/ZMo2gCjTYe4keURBWKLoge/hH0RX/b5+DIPr3mCEUHyjRAj5AfgazpAQvmpyBf0C/IyUWBuhFXx/Uq74gZE4JMILQ1hK4YQH9bsDtDSzwlPRu+ARig8ZL4PhOxGLqy/8HJSg/hMpL3yM4MEM/DGKG6SqPHygIJ1iKa/sw2LOlXECvQ5KyBrADTyiAplCf9YucoPkHKwOQHjAI3tOoTVuCQamkRyuD+aOvDDjBE7w8DDmFGDCIsWAKA0ADmCkhLAAHizskOzgDCdyDSqhAH7wQtZATPqivGSDBVpgBANoHFDzB6PuHQgAJ0CgWeLOCEsiFb3PAODiDJ6iEHuRBGYqwHySeDvAcJjiIqOODcjpCd6O8LMiA/zbUP5BowX94wUQxgHoSI1uKBQJQhQbIwi3MBUoAxB6EkY6AjzAsllngD/HxOOV7tMk7wULIgEIgAQooCGdoidvDBoMwvzg0CDlUj3oSM0tAA+dhAV4ghCgoAC6sBFXMBTdAAaArke44RANBms75iDIECebJDGOiED+YheSbPzSwBHnIgG1wQ1AYiUtMCTo0kGFCOXtDoVKjhH2YhRbIhVy4AD5AAVa4OCSQAwbwqI5ClIOIg3sZhoLQgH84gH/wgYOAln+YoGRZg634gH+oRFp8iN/hhN9hOhY4BC64xuWbOkNgw0/LgoPYjo24xGYMiYYENgPZNctLgX2AN3erJP9xqIIqIIcxiAMh4AIO4AIGmIWQnIAOOANwM0cQ4IJhEAUN0IADaIcD8IED0IBXGIAOuIAXgIOw6IoO6YoMLIj2y0eISLqRCBGWgAcTWEp46AhM2AEN6cCD4AJOgKsyOMJW4IVC+DRJhCyDUMhZLI9eOAgjgIixNIhPSA+ELAjpozyTs4TamoFcSAFLsITkK4HkC0RKSIQqMAZyCIRn6IFcGIJVKExtWAVmSMx9aIF9CERDMIRYaDcZqoJcoExxyAWAhIZ/aL+j+wejBJ4iUB8LuATW+MyN8MKLaB2PaJWCUMpZ6UEJPAh3IUnkw8p/UMJP28p/oAMyKJCyTMuz/If/TyCFgkhLAFET6Ku8FOiETvAyL3Oetro7t3IrGrMlL2sFPsDOx2ROMRIjFvrOf9grGZo6akxEGkArovuHXIhNW3mXCCLK8khEDuCFXEi+Vpi8NtyGLHjC56iPRwgLwigII1CEGLg9f3iER3CGP1CEfwCDENBETqSPJ0TIYrSIMPswj9hKhJxQSXRDY8wAJdwHXrCETrAf/uKvR5O/vKwkXkiBFh0CZvgHURgHvyGSvWGAAYiKRchRjuhFLZMYp5mFfcDO5bMESNzP+yqICROJZcyIR9DEz9NEiHiwBI25fzCCECiwg3iHJzWWtVxLg3jCgjhID21DM11CNEVB/OOH/1Xggn0wAR+ASXcsCFHgiPAhFhdAhfJYkKggEnJkCU4wBU7ggFv8m9HBjFyEiFmgpMgMBjvcSkhFSFBgh7E6iLBkCil9iAPdxEe4BwNtkyRNiSMoiCMYVSf8h1HVzyPgyoPczyyQh21ABn7YhiEABmOIhSeghAtYz1lIhzjFB5pMRzvFmH0ZFRdbBi8omqbYxX+or0RwVvqMhZHbBnmA1FOFCCQwkE2lEDH4h5n7h7UU05CIVQhYhSYjr0BI11gQB07YBk5ggHblBC4ggClwph14g3sFARXggwuohF0tgPab0XYAic4ZSpKQERD4HB8FntCJgpFwF/04BHZrBWr00P9VvYgAZS9+KIhvFQkI+NgMeCdogiZnCoQdiAUuYAN+5AA24IB3zQULyFd8fYM3sABcLQgY+wdZEAU6WAVx4II5kIUf8QiDZY2EhU+oQIXhGYmFfYhElCE/yIXbOsE2XNX7MtV/GEvheLU2aINu7YgjkNWZE1tv5QdkWIU8mIM5gIZQWNlBDclcsNeUgcooeIJoa8wn4APOaoVW0K88iIc6vQOkzIhFgFjzONr4eAqk7T0YKzpo6RxmmAVmOARDoNgUOEYzDdPFBdeCaANk+FxkQMF9GIJtcFMuiNx9cFOKtAReCMRWyEa4gqtcaIXK1U6+pYRVeIV/MCs1mSYnQhb/+FQdCayEWdAGXhAHXpCDSjoEEqWEzzLGLLDaVx1T3dzcf2iDh+haCGiDjy0IfpCHfaC8Fq1L8q3LSnJREd2HinzdQ1gFGXUAUegCs7LekXCAjNnAgmCA0FkFfphVfjhBFRomrtTQ/eRciIiurTWISzU0rDUIZPhag4CAf5DggvhYC7Zgfuhaz91gsw3bDIBLS9iGV3gF+R0HB3CAV2BNbUqDbDo3TpADPGgEGaaaf3CvEcgBwFOBaaJKNmDR1q3LfcjgUi3V6P00JwRTg+jWfBDX+YiAjLWI7mjSf8hWqMDej/BKzcDiCL5gCECGNphVYGDdyZUDBZBfs6rTf2gV/1BKDT7lCBBoHcQ1D9IgDTkjiWiCCN0THyW4AQrIyEN4Vl6INkFuvkpiXUsAsf5dBe7t2s8lYqxl4osIgbGqVAlRyIwYKyFQjCsmgV6ALAggAQp+iFBWj1BeBVlNgZ/lgljoARh4AjfgAs3skd39B90lFkKEIpRoYaa7BkAgB/r8Mhc1OXlg00/+5FUAZWS+4JnrWlR9CCRG4gzZDirGDE4GBToABRIggf78ByzWYr7AYvf9hyuY1UMIBDx4g3MGgR5QNHuslX8Y2oJYWt9VPGZ1oNWCCAEQB2i4gm04AjH4WGQuCG++iM/tXBJogyPo51EthFJllwTGCWumAyjYzf9kxIiB5ohRRltQeIU5WAUEEAcCMAYB2IWR9gWSfhGH/Qd79BH6faLJKAgYeQNjwIEryANsLmavHOhsXoV+XoVQwAEboIBwqEQKuIEbcIJtQOpCWOphkuUioeC/5aWOvd7UgAKJpoN4wGo6uOY8WAV+3gaNfAYleJEA8AUBIAcCkIO0Xmu1viiSviiPWFqYJjhCxINdeE+LIM1/QIGqUCS9/odnKIiVvsfCgBEUgJFAcAKvvoJwkAJnaAYpttR/qICiMAiC0Ay80AhYOIgC9AgIAIUECIVV+IBAoIDCNOXu5QgsruiR+NtVeKcosIBAAAEQEIAAqBqP8YQHKQg5KIj/3f5rjQidkOhtvjkdVnhpkBidMzAIvE4LixjswRaf3X6IhKABciCHZyCEKjBqYaiAc1BIZ9CJh1iBzMjsgsCLGqAHeri+giBvjMABCiDMhp7qjfVWZOjizyUBcXgRGsADs/6HKCBdm05miMDmgkhG1q7oi34IBYcsULBmXxKkALhtjwDug1DNj7jlh+gb4IkGh7AajbgXGFGCf8BroBgwRqqaSHCvjLCoXagKDAiHJNCDCmgGnfBuetjsQXgIguiHfrjsj9jx8/6HdTiHc/gBnTgHsoMIG/+BsasAPcAL9y6Iy94FJagCCsCBbcgDCf5aK87ef8gDcUCBkv4HATDp/+WmJmp6BjYnBAIQh21AAKT2gG3gZxwQB0mgAALAAnEQBydIgHgIdKwOdEGngzywaZvGZv4tBHHAAhTAss0lLIZQXI1oBBD3CAz4hzAwiE1fiqdAboPwBgt3FRTQAVdYgZuogPCuAONIAnqogRWgBlSHcoNYh4MQ8lvPC2EwO0t8CPFe8n8A9otYRiWP8n+YcoPAgk0nBKPGARwoQESX4F2KYGToajI4bCv/hzQ/2r7+iKiyCJe7AdOZ7TiOBCxjcacwCEhnuroB3pBQTRqgBYt6iE6vA5zQF4dwd6hAjMFQiPpY93/AAFfIBFo3u+sYBBrfDvHGiIUnu4X/B/Emdv+LOAdiX8bHDvaCAO9/iOyMwMeDuIFwsAEMoIGyLgZfCIAXGYNd8AVfIHF+R4iT/wcS7/SDIIeKCgOBoHKIWG4S3+uFaAiOgPRiAPiHyPksQ8+QqAVIr6AKogHFHTTMeApAQHf/6JjQ0AEMuIsVMAPtMIhLtOSvDPuHsGSd4HiLuMSsaFKJ34hwMAyQ8PiCqAhaqIWKOIhuNwiJsPmah4himPuMuAEMEAJ/H4x/mIy613eLcHpKvwggN3pF0tJZGbS6KQirZ4mrMAgduPz6qApEEIQbcAV6AA6wD42H7wiwT4Jpvgol6HmcqPuLuHuWoPkAeYrFrxDYz4iHtgjI95D/jXCWryCswEkU14eIh0wJXe4Iq1cFJIgJ4vAPW4cISx595TBvg+imlyfvTMf+hwD1gjB8g7CoedcIxIeKsKygDYF6zeB1kIiXZnsUZUF6RSEPdEiFunlpyPgHeY8POPAMOACITez6ucr071+NgwoXMlSop+HBChAnUqy4cF3FbuGkWKyILhs6htl+/TuBKELHhtlopWxJMYIUlJBc0qxp8ybOg6wUoszp8+dLoEKH3mxQcw0PG07+/LPxz5WZbisUJiRqtSNGhSsGCePosufVsAtTiaWILmTZtBZxLTyl9q1FHi3dui3LDS3cg0bXVNykUFFTM1H/JWnYrWFhi8LS/9Jb/I8eQ2GLE4djl6/XP0b/Dv9b7PWfxJq68pK2ya10SrJW3eJi+++dnZZG76GuuHNhNNe1d9P81mAdGMAHlYZLUtViOEbJMDPKly8ZO3bB/4Tr1q1w4qGQ/63Y3lDYCs3O/yVTtKJbDVcICa9wRW1LzGYtR/Oub/9gnH+pfkyMwyrafQEKOCCBBRYIxD8AHCRAfgY6+OCAAUA4IYUVFtggQx1YuCGHOUkYCU7coHAQgh2aeCKFCqK4IostuvgijDHKeBMbM9p4Y1reHCQhjj36+COQQQo5ZIUWQGTKQTUSuWRFRgnlRVm0UZQGhgIcBGIDfP2zBgVMqsWFl2GKmf8WHCD+EwAmyogFBxxp0PICC//EwsKcUagQRRQ9jDBCID0EctAYv/yyixzQKDCHQgqMuSijjRKIiRZXBXJGIIG8sQMA1Sg0iUIKKsgpp51igskUKvQQCy9+sAENop6Y6WhHYAoJwlsMCBgAILAaiApFh/xDSS4wjKCMp50qBOVByLoU6j/VAEHnP5eq8M8SJk6gK7Y0WZntUG7UElYuI0yBmrLNHgQDH9VWO+EA3KJ4bU06uguhG5do+Y+8PpVzkKakLQPRvv+oEcs/I/RowrwJK3xVAv8gqpCsC/Wb0jEpKVsuRP9OvNC0/1ygkBssvnJQFws3eq/JaimZF5Qt/4P/8csH/VvxQg8kG3BDi5g4cspiNtIzXKtw8sG4/7Y0ccVQ0myRpuVMsrFCTU+iccYL7dBiFyUDvXVLKMfo9T8a3sRBKNBw4kYRCuFMUaheTAKAlVO//PQ/y9C9kNtQ88tszActbZEyseQS5rWz/AMv12PulTATs7jwgQVeQKn3RJO4fczbAmxrLuXVgNq52gxRPhEAOxCx8pKzcJA46xaC7RMLfNtkt6YAHGO32w1NnDdFMNcd+tqh197DNv9wkjoH1yLeOlwqNvQq82nYJK+OHf+j5lB33x36pv/IDjD4B+0bfNPe/xOFOGxwcDzzQOfb/oBTxBLLFMjavKz4Xvx7//8/FSuo6cSW0TKjUYSAC/mX08Q3iYrtC3N6e4M41vcPF8DvJu1aEiBe5xLpVfAnX5CTQrDXEgkog2/3oxvc/rG5mJUDWcGDiORqsi8B7ut7q1sSAjpYHx7psCYC0JMI/8G/iVztH8YIGJRsZrSp0Q0TfNuY7xgiuYr9CxMHAQAWE+Q5hhRrc5r7x+CElMMeegl6L+KgS36WIBXEoog2mcIkxhdFoaDQSl8UgIQCwKOf8TEb/wAEILLRCD8CohGA9AUBXKCzD9yGjI6EHxpbAggJWYAFKnhhSsZlszmK5QFeUMYxWmgTM1HJF3JYhM7UsrxHshJHjXRJABRkMExWJP8YM0jWy2h5lQcYkCEE5B+UlrGv2n3xIGe4IE3K0MqU8XCZ/wBQANiIE4MxpBy9rM/9HjDEhjjvDYfgBAVm0hIm/EMGzuQWDyOBoVYCCASxsF5LOjauYAoxL9ckSg+4QIBztohX94HDjhSyTobIwJxc80NDvjXLf5RDTeNyyRB1WRZleGGbHcHZ2pRBBAKQ5Ea2gh8q5uBPR0WyIVaMUUlbMoUHUPN6LgnY/uqWTTWVw6I1M+C+pqDTmthsm7HYJ5BuyLwEmIOkQWJLKvLkxpawFCj0PIgK+MCCh760YOIKoQwVogJCnKBHHEhl+0IKq5T+iKoQbSlOHlANFVVjBLH/MIQhjii+lowADWgwWIkyyUUAWMATC3ASRbjxghMJlZ+GpUk9aEIEoZQDrVkNmADeMIVgUBYNhjBrTyfS2GCgoRPBKEdOhbg2qlKVpubDRBR0AFiGaImsh82WGhemwbSsVAVqOEgQGZJbhbCAmo3lw0HsSoWHqslmJVKDWaeAhn/AlRLIHcEMpgDaq+oWqzF7Ggho0IDVQiQQ6xqTBl4Lv8QeZLYLUcU/YoOTcdUUtxWhJv/eOoJ9zcAQwf0HMCzhWIZOgQ/zhYhd9RsIuEp3CobQbznG5VCX5lWIk6CVecUrYSHNtl3IVMhD1eCIf2w4JQgyazUPYgyGik8NrQgG/zWDcRBDoEESTajCVcelhQdMYQSGCITngmffIQCDxfYNBB9SkILlSjRZXtgBCtZglCVPuMlDmu0ExHaQSf3jw//QwhQipVeKNPYft3hGIBL8ADXcUsUKWS4VxNEEcjThGbh9QDl2MINgXFZzNravXYExBElUARh2DUQwgiAJ/IbZIpucAgrgoORFb3e7EXYypFFEA4j4YQKV/geYsBBG5E7BETutCPZK2xA3DkGuLIXrP9CMhipQYQi36EMf2vxQGt8SDcHYQSDeGlwqSEISt/iDJAzwjyr8gwop+AcYhnBLi4xvB89AwRhoQANf+KIYI1rAoyMdae5WaA+84AUlKv/RiifEYgZ7aggQVLCE2wJlXFUYA6xvodMptKIhaBhCIf7RhCaM4cvim2yql1tX5tpVEmA4iCT+AGxioyEFf7iFQti9YU9rucGmetsV3egLbXO8SScqAbhvud+GzGAGkdKyS1/6gBFDHNZVeEaNl3vmXjfhICFowi/G8KcHBGLZ96XCsP9RiD845R+SUIQkhlAFYg86BBC3L0MMsa8HNDgH/9gBiP8xooU0uOMcz7aDZsEL4FpkCXwYFxCyvpANIzfEC+lDN26B4gEH3ABkcHUfABUDO4whCjqt98/RQAUDuJohfXD6oGnu5VsMeiG80G/Wd2BjnxesvAoBqNdro7X/zA9lAt82d4YZcgj6HeTkEBlzzRgC8YPEPRhVELyembIQdywAHDzQhRL+JPPlvh4YZCDDLVYPa1g7wxljGMJBVu/lYXP2H7xIAYptFqm065QPVKDzQdzcUc6jBh5h4XaTEXqQCVyrBbkgO0PWbLDbwrMl4iDPQTQDGDBMR98H6cMoxrB3O9gBG+4whn29HtDtma8pxPD1gf7xQL/9g+zpWx/8Qs0NmwGkABXMgIZx2EG0grkZAhVY1rC5A/eFIEPkyopcC5g8wRSwwAXkQrWg3C8YA7sRDIlVhCGo2DOQQEPkQR50BC58wxr4gjj0GcIVIEMkg0JAQTz8wzxAARRA/8QYhMNBHBsVXJ+4qIGWnZ8xdEIHDtvGgZ8Ift0/xFaAeCFDmGALtIB/FcwU5EAnUMIIjFh6jYEx/AlzdcLaQcTq5cM8KMQqpIQusAX/tYYugMMYjIFCgGBD5END4CBEOEHSGZ0BAJ24aJJC0NmB8UIu7MIvqMIv2AEP2AHYDUl4+cAX7oaTiKGAkGEZJsK0kFm9/QkHMkQV1BjZ3VhFENtP2AEu6AIPxMAmuEPeAQUC6lsTkIEBLFd0Yd2f2CEwDFcgjMufvOHiyYWujGIp1sYp/oMZTUgL2AoXdMBUzQAl8MGAWUKxNUTNuRkV2FcudIJjjcsOBMMYuIM7hMP71f8EW+CCHcSAIbpDN4zCT/RDCPxDHyzAGFSBJEjiFCjDDCwXGgBDCkQi0CmEMbieO4QikRzANWIjHBTShKjGQShTC8iKVHXC46UAL2TA800gMDTeQpjZP9ghcwnMP2TZQ43AM/hCoPwD5v1DDPwDOBwEf0CEevViDNxeQ+hGQ9ABRPQiL9JHQhbMnwzOFGbAORYbFVSBOIiDOyjaP5AXrITXRqZMCxwELyzBCKjBbRlCEAibAQDDRLwYnzFEEFiCZ43LxI0AIbiZT/4EgBzEX/oEK3zDP5BBMwacHQbBP0jhFAKDnlXB9i3OWE5mgTAAGqoBNRkCMLTlQihmRUzk4Fn/JRgZgrlV4jOQw0L84YA0wRUMARV4pkLIgxhkQQaopAE8Qxw0AG2AJUZSpm+GRSX8AwMkwghYQcF0giUIG0V4JgQoxEQuRK8tRC4Ywp5MlvYF5YCAg8G55kIYQAZQIFxeljHswnaBpeX9JnryBhfwgQXG5Fu+JX79A2xWRAQyBCIiH8IBQxXkQhMEAjio14Ak3WsexBBkQBAoJtAFg/ygQKMxBGCpQtr8yB78w4SmJ9AUgPOhpRocmAG8HzDA53x2xBVcgdFJgi8sAD/+wyiAwyDGwNZRo4AM5EEAHTDIg2MqhJ+JizEkGbc96G5ZKJAKRXCGyy21JXy+3/u5ZEvg/+K+bYIn6gKU8gArvBJ9EEWV1kS+HcR3hmiqiUss8KjXrJaRBEmFBql9NBOB9EAGlgEljB1mdkIKfOhCwGVOFI9O6AIrXKlSBkgwpkAW/INyPmeCeimDZklO9KSZJupEMEErXEALuKHBJKc4xOk/eChQGGJF7OlN4OlVKOZhzmiXTkEuKIGSbddChCKiKmrroOmAPME/NCoamptJvied5sTgVQSnhsUrdQSAMgRoHkSgBkEwPGMuCEKpqmJFpKqqLisT8EGbmhsffFskVoFiCpuSuoRicmmF1OpEICiKiSo53EOjgZ84KQTKLSu6MoQMtil0mSQvUIGNLaY4dCi3UP+hqNaBuJpquu7rTajAHfBCJYxAK1hCCgzOCADdW26hct7HrvLGFKKYGjxBuI6rQgAWJKgpuirDj0KIMrWOqybC2M0AckLdwfLCWx4bfhnAwnLrkkgkxPKBJ9hBluhrK4kl15RBx7YOE3ybf7VCve3JDEgrkqIsrLzmXU3BDDwDD1CsYY2DgERohShTGQzW1owIHzzBo5acuZXmLU0qXMLlBAKqW1oEnUaifBoIy9bE0bKAMfxCA9RDgzJEuSqEcSZOOwwIp3DSsj5BK2St1oqcIURkRDYE0TKES8JlENzoQgCdOdYqXF4rUPAAZ+AXXAJdtmprR+RoqcSCEByrk9z/y9yWQPdMSI1cGLb8Db/+AwjECdZSgtYuQWm2gpANrk1MJJ0CgzhQwA3s7kFQAAVgwFSYAVEgARR2ptkeRFsmr0VwaY9VIQs8gy6MK2Ahq4OsDJIozPekbt+67t8aDJxO4LEt7ESIL8JtJQZsgjM0w0OkxWGww0GIA5/xmWNu5kGkrU3cJWYSgipI75bwBMn9w0lBSOmmLtCIrt+WQcnRCZzO7mJ2xLE5JgXQXm5Mgz+o7/qqRfFmwgq0hyvgABmIQ7b+hDkyVyCkpRsoARzwr0LUxYmwD5CGzKuyThpQLRM8arkhcAncEiV8p5C5BO4+Qww8Ql38gB5cMG+kBxkk/yfy5oRiWgK8BsLAPIPbqvA/sDABV8jHtE4Z7GzIIvCyLfAQEC35MsQDh8Mo4MI7vIMFB0gN3IA4JGetYm5KHOieYKYxKIH0AtZOBCdEkGB6om7qlgDIsicCs2dMfmcYi+ZCFC5DAEMT/IAaF7ERMwQs5EUbi4Pjnq1NfG2XqkEOlAAhgEMe64RQcMQ0IEKkFUtplOWEVUsJtCl75jAOLzAit8SHAsMNaIL6ekd96EEzrMAHG51VCGuN5UAuBILnOgkunEEY5YQVXzH3zcAFYCIL5DAhd8J3ZrNLHJs4EIImgMePIK47puUMGEME5HEDLPNCXEAW4wTVQvNEFFZFuP8q/EiANYMbCyAwAsekkGlzSjCyDUzFffAANRpi0Q0FXEKsWz1DCkvvMjfzQuBB/9rEAMgCPDfE9fLTn5RBtTxrIZec7NZmgRboPygyiqjGT3ZqMGDmCOQCCvjGuOrCC2DoQfDxRQ+F4TTZEiwBE3jbDOSwNUerSJv0ingHSP4EfAKqJASBuWFmLPxVTCsBTaPrPRlImbLOd/WtBs4Ae94SwdZmBuCniwgDf/gDUYytAXSCBUJXLkzxdoFDIBTAhO4BRC8EjDYEFtDE3crzTTtSx5ZB1lqB1vIzWCMfUbfET/rDUPqIAdjlnixBK+TCCehmA+gCChTABVRCZrdzX1v/aBmI7isnQixrrSGkpEiX9J8uxAJYBH/8QAwsNpAIK0sTgHZV9mVvtk13NrdwNoWILldjIuzOAAKjQUqmQG1mASOz9j9EQErDdo94qCVArDiSwxrEwW1rNjtTAgwwBFhUBCB8EEXcrW7jNGmI7oTWNYU8aw6XXDBgM1hnQBaQAC7WxF13Bn9o6k34Q12YtX0ImyXc1Z4cQhX4AgrkQi5odiUcOAygQG4eRE+s0ngTiASUhc/l9oQoU8hstRfDKVhnQWqPgTOEBS6YZ0uU69zuxtgiL4rNAAscgoFndiUgOAyAQBo0WgTIgXBe4zJ0XWnwtViYblhUKHqHBTw4QE4Y/xQMcAEvlJwXB1mHZwEdkIFVYMM/UPk73MgEooG5xcIF7EMLJEJm70ElLHhubpcUIJQ3spZCXMJBWPQ/iDdFUG8psvJBgNUbwQ8LfJvrrvcMfDV8pwAO+sVQUHlF8MBRr8iQbS0lGA4vXMATMAEINHQDSMEAcAEDVPoEcMEA+MEZ6EUaCMAHyYIGjMMBhJdYindw0oCy4sZBSINVaMDd2mwFUZBNWHj7JAIXcEG5cXV9mbaHH8FBbF9amHV9I/pietYI8IG7psAhEIIvxIGSCUGu5zoDTMAsbDqpbtenfwECyIIowLoGHIAPHMA4aADCeAxPKhlE1IN8RDjrHAIvcP/BOPI6cYc1cmcBidZESt8ED2DnvvP3T6Z0vzelQhA6QxiEWIg18qXAf0NXK3ybJeSCi1cBIVC7pU9AtfuBDpTqtnOBt5eCBmiAD4R8uc/BACQ4jzLtP4AfknyURVz1QrSDrDvZ4Nj6TYyUCZz7TSzViewTB/CCBm61IRw3vhXCDq42XHR3QyjCJxhBcCiCIgSH8B7EJyAbYFT90ovFsRHt1jufAdRgslPCo/IBHxx4C/DCLHDBLLRABkQBOuhCHDRCALzBNqSDLMTDMMxD3g9DOqTDKgxBmwILISxdm+1lGASCL+jAALj8BE3ENTQK1NqHj6OGztMEeL8IA8yCOAj/t9amJG3SJjI0zGqv9mfkhXRQ/UIYAeo3BNbvhlgvsvNVoC21ISW0gn/tyQig5Qj0lp78Ax+UWy5cgO2zJ9kDF9m11O7HSZwoRLwriQsvDI+jBgxXRHDaPE6cuwl4X0f0wEm9gULIIFFkb1kwABfsQ+3zei6Y9hF4OATkASLaR+tPRPyvfoD8qVXevyXUoC29bnECxAg1A9VMIahG4AwrM0bMmMHnH8QZ/2KN+Pdv4kWIF/+NKMHHEi9mHLT9k3YxDsd/KlS2dPkSZkyZM2nWjAnEgk2dO3n29PkTqEsv/4YG3cmr1cMZnXjty5Ali7whRqm6NPLJyL9P/xR1BQOG/xRWrRe3bq36curLDDMzGAiCJukIuXINThE4wu5cNIaoBDFg6R+vFIIJD7aEJljEljNYOGyVS9wzFMV2vXnTMWIsldDOdvbcEshn0aNJVx1aVEDpi1xm8XrIpxWlDE+jZlG9E5sdHthCXFT0zxa2b/++YRsD5lNZMN3s/Lj9c22GFIMNULHUKlgruJaCdA/MMW2GtFlmPy1PPgMvS51aYXTv0KGhTpRyHSqQ68IFijNKXFg17LkAaQpNwKr0KxDBBFdjjRI+HupkNqgKyaIQBV3ChaNH/vlDpW4e8eedf94pbp1u1sHGQpue4ki6qVIwwABgYnQpPJdsy2IIHHWcbf+I8qbjxQBDDGnFEPiMmSGWGYLhgxJeMpCHH37oiKclDVJMkQGVJjjLFI66vBLMMF3igBcHHXSSPHmy2OYfEv7pYwGb4vwpxJgeeWQdMDhSZAwM63wkRH8wvGhQMWlKyyfbbMzRPB/L63G2FIZIwdHZoNwmHSv/8eEfDUQZx6Yuu9wgQTw+G+CsLP9ZZFVDXQ1zllkSUaqTFNKMSh6efvlJwzpjyi0EPRX5JLhXLVxLURv/2ZG8ZhvtEVrxxFuTH15y4SWdeTTQwAcrRflnFZk4uMgUUhO8bDRVq/ryH3aNfTdALli7wMFWeLkVqovoCIejOV2K019/bfJVpV7/uRP/mxg2cYaHewiGN8Fcj1AWKqjMcxbH2cTgh5kULHnigicKaCGdYbbF56JvOZnJXVLngHgndWMqiiZWgToQ5pxlGoCLCbiwNhY+OulxQglV2lWmGBaIQTVcNAQUpkJ1nli0XK1m84htjpAna362iRKZKOXhQhxgRggEABX6uwC/AmaRRRRNQe1UJxeu/ELnnnDGOW+eAhBwo5ZmmcBnLoI2hGgKb4wpgpaY/icCpS30R8S+L6LaqMX/CbsNedITxw9toFlFm1C2CYUTTnIJZIfWW7cAExVkwA+/SjiA2/Lcf1JDd54wkWmZB0Tj+yUVDskFNkuezHHNf3J9yRmZpEhQ/0PKexfjH+x/WnMVCLgwZoQ3dqjG9Tu4SJ0BTjhYhAEGDlEBkx3Et6wItfOjnY1/uvj0H1FEKaULNEFAZ9DVOwMaqwgXEd4/JpGaqoDsIixwiR8S0YF/JOIQDrIEpYxQMee9RGCvsl7ftIcMMbThcjpZCwRA8Y9b7CIQbwjEFFjHuh0YQ17qUx8H2vcBC7QufuL7guxClp9EXMQBoohHHkLxilf8gwA6cRdPCnhAKxrQHP9ARVVQ9Y9Z/OMDRCgSJWzFvHypZBRX7BsyeFKIifFjFfw4gjhiEYgYvs58CGAfB/jYPjfAbgdfCOQbvmCBEkTkAvaCBh22MYROGIIXr/+IRwJ2Mi4LgUCNmRSQArb4E5bApANuOAQlluIk5qmJTZq0HAp3coQj8EMlR7gCBC6CjG1cIVza4ET6+siAP85vBxepxj9Y0KR9tKAF9OKDIfiQC0w5wCcyU+U0X0JJavpkS4nIBRFysRRK0SZZ17zmKyEAARKsYhXI6F4c50gAQuAAAe1jRpZmYTjWTUEFsXgCL/hJHz7885+taEUnOsGFOcQDmlHYyRTFeREHGrAUHIFmQznyhIsw4R8XOGQi1MWFf3iUF4aDjQEutiKKjjN7bTDnPxo5BF6IIxfXYsY2NsAG0mkDp7xoQT8pcQH2CLQVsBGqQHMxBEk6oAseOGn/UB76j0boLoAXiepSL1KJSsjgIlviSKyY0aDkRehiVD0g5mDSBn4gYzbqsU5Mc2EJtuZioPOJzVwpMVCgBhWvfBjCy/4R0W1UUayBVYkJptpQGFj0Ai2Axiz24cWPDgGmuSCoISjlOQ/eyKSCnRpHnteSNrQBGSqlJT+GsA/1WGI9lOhELgwhWbgOiT2unQ9BYYOtV0DTAU90SVM1GxPe6myivc2oDC4gEvXwE7VNctKT5LGN2pDnIlCRR2dBKFyIkXVzEEAGBM66XViKzXPhnW5z5SGG6e5jHwTNxSxWEY8uINUBJvgH3qxbX3FKEAYqUUYumAENBmzja1ESsBgM/zCVXDXLYjIZwz+QcJHoNc6+FhKD9i5CS1pmV6Wi5S53kXGECXdYDK905dbW0wlxbMOJXXiv/i4CgAgvFR4sFmt+L6IMjpxYG/x4EWpzQQVgONeyFzujS6pwkQaDCcIv5ghoOWLhckJAw/wA7ZRDe9aNZcEA/yjqHF7RhS6vWMk9gcM/0hBmBNHAqY2IBEdM9Y8cvEQO/0gdci1BCdVy7QhZyDOCNdcSNxkrei9JsoAsHCY2VrjC2y1nhrnbBjF0OANBuNYsBqCAL+NWQS4286Zt0uaU/CMSAaAvMYnJgh70wA8cSA8vmkQJ1GbgCI4OcZ73vJZlhRNegQYTCg/95P9DI/oifxYNLX+tkgs3Gcob5keurMMMXjyBCHNIgJdbwgljBOgNldH0AcfM6dLY7B+X+McYMBAGFKDAAioYgT75OYsWtOa4TQoJL77GYWR0eMSKWhyu/2FrMTUuhAVCIQpZ6KZZHttQCGcjG6PEz6bkIhYwcMMAEjDtGHf5H3ngCGBFU8A3bDt3Y4ZDmXuyi4uY/CIwUDmNvd2SWjyDAsZgpkDZo1o78yIRqOUFMHpUzjhC2az4ppqacD2xCrXkyBcJOKCVTpMF94QEdHATMkhAyyvERNi3ufCxwyYOSfFiBDvIZyy26dEBcuQGLa9JmUn+k4dKMEx/y1sjAlGFIv3/c0jyqTMvnAdHOJpT0cn+7L1TuKyWGF2TFfjH0lsiBKBEnQ4trHrVxeQmYmdgG7wwhrZB0AMY3AEmhVW7S0jO9tHfJg2AiMQzeGEIS3iua/zQLgRwaU7bP5nXm2NldC9HNexeEWAxGcPTffJrNoIiH3RoEwmybqErnHMbsUABHqaPBwCAQKGgvwhf/2HNi6Dg9AVi+egB0ZJiVGEIQ/jaEe6tXZW4Cf5tasmvS0iCWbtyWfgPv58vAgpQ0EH5/C/rmo8jCPAfEG4mri7j/G8VtiEKdgEPdkEAJNDkMGn/LrBv3uDEGrD9ZonqVCJcEPAirOwf+IEE2GgbCiEFYc2N/57n98xMBFvC/wBQJVpI4/rv/V6C2Dhi4SBgFUBhDvJgDkRgG3BAHOSAAAjgAQPAFwJgF/5GAMBPJ+QOA6vwLNIOJhohNUwlEAgAl06wnCaPlsLlIq5OAdmo6kDhCpzgH5wABwrhDVOQTdjE366pCf7BBqgiBuUv/lpIX/4hH/4h8iLPD2npz84JFH4QnRpJHMQhEEDAE5JQHAgACZGQAM4AD9oM5XqCCq3wJwKgzTiiB1Ri+k5qFD2BJrpoJ1ys7rbhB/9PEYHQBsOlkQjhGbYhD8hgBaRgARZACprhH6QACTIhHG6ADG4pBQshGUgjEy4CFv7hGYGiDl2C9vIgD/9E4ApwCRS668LYaA958Czm4R9ewRohiwCqwBiiINsCgB0DINSYMAqSkAgo0ULizBNjYhNlAs2CQqne5QUuAhVLAwsuQg7kYACGYICwIBBQYBca0hf+oRCykQIq4AfO4R+cwTmcIxj/oQKiJxMoIBycoB+MzIo6TJ2YqAEbMQ+uoAODwg91AgDjoQEJ4Qxe4AUs4AXwQADYMdR6MgDOAIxeQgrvMUweCigvQqHESqH+8R8CgTSOkgIIoSVQDgWeIRuv4JYmshmiBxhfohmSQCWo4SI24VUGQSd2jwTmQAG2AQv+5hbRSfYqbPJykCpeMlwAcBsOIRCiwAJAQAIjATD/3ZEjLDAoL+IDCGEoO/E2sDDMVEEnxI3NOMIpVeK3OOID/kEqCSGKDOgoPUMxMfMlLgEFsAAHtoETbokfrsAVhKEZLFLXpuci1uEfVsBCovEfaqAmzGEbOiwmSuis/kENn6EhTU4AnkEc0AkMv5H/gq0Aa1D+/I8jQIH5FnAVIkMCeRIwJVMqq+AyOUIqqSIU6+s7f8IxdwIy26wz/0EK91HchpIoVaI78YAGHrITMYACtuAcKmArOcIiFQ8WaNMl1IEj+oEdxNIncPMiaoAe6KEC9KA1/6EZmoEeblMmBgEHBKHurgCWUqmWSmgE720VquAJ9/EfHjIKNlA6SeD5/8zp+ZjPnJgv/oATOONP2EighW4UOMNlFf4sncSBEHahFpwKJrrzIkwlPKsiPZdqPH9izWriby4hACAzJqRUJjDA2yKhEZ6KJi7hIR/y+0CyAsL0HDTyH86hBgD0JajBQM0yKPQAQrvyJX7gB/RTD+jhGdH0H1zhBhxPAJSgCjgBLuWolpbM2PJAHJ7wCfFA7lAuCqrgxFxxFURgFfIAFIQQAOnAGv+vUid1DjBV+TIu8ig1DyaVBBiBRWcPl1ZBAa7gBnxhzQaSNII0wmAVKNSsJrJTVi9CCVpC3HI1Jp5hNLTUcpr0Jx4S/JRACSggE4RB8S7yH+ihBgZhBQaBWv9pk03/oVo5wjZpYkLPAU4v4lthYit/IELpIQme0UJdQQd0FQtskQKGIBRmif1g6SW2ixEc0QmZ8BJMDiiVAPzObQLF7RmslAL+ociqoA5U4m984RkQYBs84HRCQVIn9mEBTP0akRDIoSFbIgzC4D2fo/x2wlf/gSk1q2RdBc3ALwwoIAnC1BnyswbO9D9XgGapYRAYlCMQlCZgIQnclCPI9CLIFXqAEU7hdE714Fo54hmwYCCxoAooAAf+QVJVVAHlkthAYRtEVAAugQZQYFd39R939R9+sl2/8zIxgBzW1UtVImpdom3PAOVAQFEvAktBrSao9GOpQlhpwhtaYl3/ayJhPfYiEvYiSFQmPkBwzc8lbNUb+rYz3PNV/pYQXGEdKuAcLPIimrUGXCET9LMlgFEPkiBa8fRZgxFzgzYmutIZwlUlWFdnH/JvO7YO7PMfbsB2cQAHQiHjJnVHcWkE0ekKqiAQaGAhddUlPCFxOeIMSBQygfUlovYGzgCTmFIK14xYaaIY/qEYtjdvFeQzfcIpDZcqrIFurUsHwsAVWjZzM5c2mVXx+vMlzqFOk4AefJYjRUPXylQKpvUfBOH7OPYiCrZ2bdd2KQADAuEZYE4cyOAYh8AIxeEMFnJdxfYfamFkL8Jj/Td7awIHboAAlOBkaQBvdaIYaqGEN3gm/1yhezmiAS6i7TqDFlKBFl4iYQm3KlDYqUJ2NP7WJsT3NnSgDm4gE+yXHlwhHN63JU5XJRQvfx2sTAOEdG1iM9dWe1WiGHyBBnh4XYeSgv/Bhl+CilVYjPNUPcu4jGshS/9Bh52UI653hXXi06gCBX6BFtBhJrr4LNaYNHwBcmkiZONAF0TDV8HPFVyBHoRhcwdB8ZqVI6JnkTmCkV0CNmHCIk9XiZ1YejhCGFriDGq4JQpWhQVYcVE4SKW0j/9hV8lBJfxXbFHYF/xXJs6NI8BvhnvigluCXy6CMd9Yb2Fig1NBQBwzZMuPmG/jlFWCBuJ4NHwVzdAXBwrZfnVNmv/jdya+NZIDbXoscpKdwRmQuJFr4ms5wkpVgjbH2SVogXxrAW+P+SV+IRuq+CJgOSZ4uHAvQo9vVXtrgXx52UJ8GCiieCdSIg6UmSpowKBPABF64oU7I6FPQJzNYDVjook/4xwmuiWaOH9x037RTJ4v4g51IlffGWlc4pZfoqRfwp8NpZZhhhbmkyOwuESrottejKCpInsRwaH/IaHFJBJquRaEoJAnVBg2uSdkszMsmiaatWBTmiaC1BqyYW9r+Rdy+h+ourdWmjRw2CdIdB9rAauNYqZ7JxOaUSfKkyOuIY4XGigQWiWsukDigORSYZ9PIBzSlyPWgahT5JJlIpL/fZYewoGHhcDxOGILaMKsVYF835kjRjrCdro0GuGre+KgawHNfmFvZ6LBki4mWngn1uAfWpizLyK0ScOtU0RLswEdVMGOFzuyfyKsa+IkpEGgEYECzCAJwPIfcLsmIjmSg0LXensmKheSV4CsNbsm0OEa/sGOV1uxq9q5faIRmjtA7lm4ThomYNO4ZWK0acKzWwK0G6C7X5uinvoa0GG1/6G1CwQORg4O7AADGMEVcFO3/2GT8zom3BS4r8S+ISeLYUITauIasiEbzFqnd4WxXSXJBi1vGa80uvsfxNsngBle0CGO0UHCJTxFouEf1iAGnAAMzIBfJtQljHonSPxK//Bak12itDmCLP/BrM3bvFUioSHBJ9Bhn1VDwYkyx/k5JlKhpjP8wf9hE5zgNxQhHFYgHPilG/j6fi1nvyfZJTQhu3uHGyDHylVDFah7miJgx6+IB4DiFNTIwXeihZecQ/DQDJxgBXBbxGHCxGGGxDOhkIWLByAhFWicNM6bxxMEw2eiyz2jvF38x6sCtEW7JsDAFjjCDMwAoGFivlM8QezXJcByE1aADZeRjKWAG6B8muI4zFVDz6/JelLhy/8hFShHal5iu9+F5OxAJ0p9NKr8IgKZNMZcuy/iG0ISOHzjH7oBN5ecJjbZxFHcJfY7QMhyAXrjIkiBI1bgr12BNuybgcZZFybAASX+gdZh4gd44M89Q9YTJNtvgxVoYtxFA0PKPZOqPBpw4SRgpt0t5Bts4DcUndFF99Fz9iK6wcOJ3AxsAMS74bbX4dHv/SUIftLXYayTgKiJWjaFIQmIkRGg4CJ6IRmc4Mix9VlXoJA1QQogARg5HSZ0IZDf/SU+vc/zNpCBtiVYgRvCvTM0BBc0XI1cPRog3Fhs/jlyfd59wwlu2ybCgREYYeIDMR/yoRd6gRQYgR3YQdk/Q8TtWiXquxvMwCXMIAQAHjep/h8y4UypYRc/3SZcXcniAN0D5ORVor3/wQ5wviUCAgA7 = 1'b0;

endmodule

`undef Mips_Alu_alu_Data_T

`endif
