`ifndef MIPS_MIPS_I
`define MIPS_MIPS_I

module Mips_mips
	( 
	);

endmodule

`endif
