`ifndef CONTROL_CONTROL_I
`define CONTROL_CONTROL_I

`include "../Opcode/Opcode_Source.v"
`include "../Opcode/Opcode_OpFunc.v"
`include "../Control/Control_Control.v"

module Control_control
	( `Opcode_OpFunc_T(input) opfunc
	, `Control_Control_T(output) control
	);

always @(*) begin

end

endmodule

`endif

