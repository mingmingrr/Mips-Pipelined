`include "Mips/Pipeline/MemWb/Pipeline.v"
`include "Mips/Pipeline/ExMem/Pipeline.v"

module Mips_Stage_Mem_stage
	( `Mips_Pipeline_ExMem_Pipeline_T(input) exMem
	, `Mips_Pipeline_MemWb_Pipeline_T(output) memWb
	);



endmodule
